module ROM3
(
input clk,
input [11:0] addr,
output [7:0] dout,
input cs );
reg [7:0] q;
always @(posedge clk) 
begin 
case (addr) 
	12'h0x0: q<=8'b01110101;
	12'h0x1: q<=8'b11011111;
	12'h0x2: q<=8'b10100110;
	12'h0x3: q<=8'b00111010;
	12'h0x4: q<=8'b10111100;
	12'h0x5: q<=8'b11111110;
	12'h0x6: q<=8'b10010001;
	12'h0x7: q<=8'b11000000;
	12'h0x8: q<=8'b01100011;
	12'h0x9: q<=8'b10110000;
	12'h0xa: q<=8'b00110111;
	12'h0xb: q<=8'b11001000;
	12'h0xc: q<=8'b10011000;
	12'h0xd: q<=8'b00100000;
	12'h0xe: q<=8'b01110111;
	12'h0xf: q<=8'b10101111;
	12'h0x10: q<=8'b10100000;
	12'h0x11: q<=8'b00000011;
	12'h0x12: q<=8'b00100000;
	12'h0x13: q<=8'b11010001;
	12'h0x14: q<=8'b10110000;
	12'h0x15: q<=8'b00100000;
	12'h0x16: q<=8'b00001101;
	12'h0x17: q<=8'b10101011;
	12'h0x18: q<=8'b10100010;
	12'h0x19: q<=8'b10111010;
	12'h0x1a: q<=8'b10100100;
	12'h0x1b: q<=8'b00110111;
	12'h0x1c: q<=8'b10111001;
	12'h0x1d: q<=8'b10010110;
	12'h0x1e: q<=8'b10110000;
	12'h0x1f: q<=8'b00011000;
	12'h0x20: q<=8'b01101001;
	12'h0x21: q<=8'b11101100;
	12'h0x22: q<=8'b00100000;
	12'h0x23: q<=8'b01110101;
	12'h0x24: q<=8'b11011111;
	12'h0x25: q<=8'b10100110;
	12'h0x26: q<=8'b00111010;
	12'h0x27: q<=8'b00100000;
	12'h0x28: q<=8'b11000110;
	12'h0x29: q<=8'b10110000;
	12'h0x2a: q<=8'b00100000;
	12'h0x2b: q<=8'b00001101;
	12'h0x2c: q<=8'b10101011;
	12'h0x2d: q<=8'b10100010;
	12'h0x2e: q<=8'b11001100;
	12'h0x2f: q<=8'b10100100;
	12'h0x30: q<=8'b00110111;
	12'h0x31: q<=8'b10111001;
	12'h0x32: q<=8'b10010110;
	12'h0x33: q<=8'b10110000;
	12'h0x34: q<=8'b00011000;
	12'h0x35: q<=8'b01101001;
	12'h0x36: q<=8'b00000000;
	12'h0x37: q<=8'b00100000;
	12'h0x38: q<=8'b01110101;
	12'h0x39: q<=8'b11011111;
	12'h0x3a: q<=8'b10100110;
	12'h0x3b: q<=8'b00111010;
	12'h0x3c: q<=8'b10111101;
	12'h0x3d: q<=8'b11111110;
	12'h0x3e: q<=8'b10010001;
	12'h0x3f: q<=8'b00100000;
	12'h0x40: q<=8'b11100001;
	12'h0x41: q<=8'b11000100;
	12'h0x42: q<=8'b11000110;
	12'h0x43: q<=8'b00111010;
	12'h0x44: q<=8'b11000110;
	12'h0x45: q<=8'b00110111;
	12'h0x46: q<=8'b00010000;
	12'h0x47: q<=8'b10100001;
	12'h0x48: q<=8'b10101001;
	12'h0x49: q<=8'b00000000;
	12'h0x4a: q<=8'b10000101;
	12'h0x4b: q<=8'b01110011;
	12'h0x4c: q<=8'b00100000;
	12'h0x4d: q<=8'b00001101;
	12'h0x4e: q<=8'b10101011;
	12'h0x4f: q<=8'b10100010;
	12'h0x50: q<=8'b00011100;
	12'h0x51: q<=8'b00100000;
	12'h0x52: q<=8'b00010100;
	12'h0x53: q<=8'b10101011;
	12'h0x54: q<=8'b10101001;
	12'h0x55: q<=8'b00000100;
	12'h0x56: q<=8'b10100000;
	12'h0x57: q<=8'b00000001;
	12'h0x58: q<=8'b00100000;
	12'h0x59: q<=8'b10110001;
	12'h0x5a: q<=8'b11011111;
	12'h0x5b: q<=8'b10100000;
	12'h0x5c: q<=8'b00000000;
	12'h0x5d: q<=8'b00100000;
	12'h0x5e: q<=8'b11010001;
	12'h0x5f: q<=8'b10110000;
	12'h0x60: q<=8'b00100000;
	12'h0x61: q<=8'b00001101;
	12'h0x62: q<=8'b10101011;
	12'h0x63: q<=8'b10100010;
	12'h0x64: q<=8'b10111000;
	12'h0x65: q<=8'b00100000;
	12'h0x66: q<=8'b10101011;
	12'h0x67: q<=8'b10110000;
	12'h0x68: q<=8'b00111000;
	12'h0x69: q<=8'b11100101;
	12'h0x6a: q<=8'b01111011;
	12'h0x6b: q<=8'b10101000;
	12'h0x6c: q<=8'b10111001;
	12'h0x6d: q<=8'b10010110;
	12'h0x6e: q<=8'b10110000;
	12'h0x6f: q<=8'b00111000;
	12'h0x70: q<=8'b11101001;
	12'h0x71: q<=8'b00010110;
	12'h0x72: q<=8'b00100000;
	12'h0x73: q<=8'b01110101;
	12'h0x74: q<=8'b11011111;
	12'h0x75: q<=8'b10101001;
	12'h0x76: q<=8'b11100000;
	12'h0x77: q<=8'b10000101;
	12'h0x78: q<=8'b01110011;
	12'h0x79: q<=8'b10100010;
	12'h0x7a: q<=8'b00000000;
	12'h0x7b: q<=8'b10000110;
	12'h0x7c: q<=8'b00111000;
	12'h0x7d: q<=8'b10100000;
	12'h0x7e: q<=8'b00000011;
	12'h0x7f: q<=8'b10000100;
	12'h0x80: q<=8'b00110111;
	12'h0x81: q<=8'b10100100;
	12'h0x82: q<=8'b00111000;
	12'h0x83: q<=8'b10111001;
	12'h0x84: q<=8'b10100011;
	12'h0x85: q<=8'b10110000;
	12'h0x86: q<=8'b10101010;
	12'h0x87: q<=8'b11001000;
	12'h0x88: q<=8'b10111001;
	12'h0x89: q<=8'b10100011;
	12'h0x8a: q<=8'b10110000;
	12'h0x8b: q<=8'b11001000;
	12'h0x8c: q<=8'b10000100;
	12'h0x8d: q<=8'b00111000;
	12'h0x8e: q<=8'b00100000;
	12'h0x8f: q<=8'b01110101;
	12'h0x90: q<=8'b11011111;
	12'h0x91: q<=8'b11000110;
	12'h0x92: q<=8'b00110111;
	12'h0x93: q<=8'b00010000;
	12'h0x94: q<=8'b11101100;
	12'h0x95: q<=8'b01100000;
	12'h0x96: q<=8'b10111110;
	12'h0x97: q<=8'b11100011;
	12'h0x98: q<=8'b00001001;
	12'h0x99: q<=8'b00110000;
	12'h0x9a: q<=8'b01011000;
	12'h0x9b: q<=8'b00010100;
	12'h0x9c: q<=8'b00001100;
	12'h0x9d: q<=8'b00001110;
	12'h0x9e: q<=8'b00010110;
	12'h0x9f: q<=8'b00011000;
	12'h0xa0: q<=8'b00011110;
	12'h0xa1: q<=8'b00100000;
	12'h0xa2: q<=8'b00011010;
	12'h0xa3: q<=8'b00000000;
	12'h0xa4: q<=8'b00100110;
	12'h0xa5: q<=8'b00101000;
	12'h0xa6: q<=8'b00000000;
	12'h0xa7: q<=8'b00000000;
	12'h0xa8: q<=8'b11011010;
	12'h0xa9: q<=8'b11011000;
	12'h0xaa: q<=8'b00000000;
	12'h0xab: q<=8'b10101101;
	12'h0xac: q<=8'b00000000;
	12'h0xad: q<=8'b00000010;
	12'h0xae: q<=8'b00100000;
	12'h0xaf: q<=8'b11001110;
	12'h0xb0: q<=8'b10101101;
	12'h0xb1: q<=8'b10101000;
	12'h0xb2: q<=8'b00010000;
	12'h0xb3: q<=8'b00000101;
	12'h0xb4: q<=8'b10101001;
	12'h0xb5: q<=8'b00000000;
	12'h0xb6: q<=8'b10111000;
	12'h0xb7: q<=8'b01010000;
	12'h0xb8: q<=8'b00001000;
	12'h0xb9: q<=8'b11001101;
	12'h0xba: q<=8'b00100111;
	12'h0xbb: q<=8'b00000001;
	12'h0xbc: q<=8'b10010000;
	12'h0xbd: q<=8'b00000011;
	12'h0xbe: q<=8'b10101101;
	12'h0xbf: q<=8'b00100111;
	12'h0xc0: q<=8'b00000001;
	12'h0xc1: q<=8'b10001101;
	12'h0xc2: q<=8'b00000000;
	12'h0xc3: q<=8'b00000010;
	12'h0xc4: q<=8'b10101000;
	12'h0xc5: q<=8'b01100000;
	12'h0xc6: q<=8'b10001010;
	12'h0xc7: q<=8'b00100000;
	12'h0xc8: q<=8'b10110101;
	12'h0xc9: q<=8'b10010001;
	12'h0xca: q<=8'b10101001;
	12'h0xcb: q<=8'b00101001;
	12'h0xcc: q<=8'b10100000;
	12'h0xcd: q<=8'b00000011;
	12'h0xce: q<=8'b01001100;
	12'h0xcf: q<=8'b10110001;
	12'h0xd0: q<=8'b11011111;
	12'h0xd1: q<=8'b11000100;
	12'h0xd2: q<=8'b10011110;
	12'h0xd3: q<=8'b11110000;
	12'h0xd4: q<=8'b00000111;
	12'h0xd5: q<=8'b10000100;
	12'h0xd6: q<=8'b10011110;
	12'h0xd7: q<=8'b10101001;
	12'h0xd8: q<=8'b00001000;
	12'h0xd9: q<=8'b01001100;
	12'h0xda: q<=8'b01001100;
	12'h0xdb: q<=8'b11011111;
	12'h0xdc: q<=8'b01100000;
	12'h0xdd: q<=8'b11000101;
	12'h0xde: q<=8'b01110010;
	12'h0xdf: q<=8'b11110000;
	12'h0xe0: q<=8'b00000101;
	12'h0xe1: q<=8'b10000101;
	12'h0xe2: q<=8'b01110010;
	12'h0xe3: q<=8'b01001100;
	12'h0xe4: q<=8'b01101010;
	12'h0xe5: q<=8'b11011111;
	12'h0xe6: q<=8'b01100000;
	12'h0xe7: q<=8'b10101001;
	12'h0xe8: q<=8'b00001010;
	12'h0xe9: q<=8'b10000101;
	12'h0xea: q<=8'b00000000;
	12'h0xeb: q<=8'b10101001;
	12'h0xec: q<=8'b00000000;
	12'h0xed: q<=8'b10000101;
	12'h0xee: q<=8'b00000010;
	12'h0xef: q<=8'b10101001;
	12'h0xf0: q<=8'b11011111;
	12'h0xf1: q<=8'b10000101;
	12'h0xf2: q<=8'b00000100;
	12'h0xf3: q<=8'b10101001;
	12'h0xf4: q<=8'b00010010;
	12'h0xf5: q<=8'b10000101;
	12'h0xf6: q<=8'b00000001;
	12'h0xf7: q<=8'b10101001;
	12'h0xf8: q<=8'b00011001;
	12'h0xf9: q<=8'b10001101;
	12'h0xfa: q<=8'b01001110;
	12'h0xfb: q<=8'b00000001;
	12'h0xfc: q<=8'b10101001;
	12'h0xfd: q<=8'b00011000;
	12'h0xfe: q<=8'b10001101;
	12'h0xff: q<=8'b01001101;
	12'h0x100: q<=8'b00000001;
	12'h0x101: q<=8'b01100000;
	12'h0x102: q<=8'b10101001;
	12'h0x103: q<=8'b00110100;
	12'h0x104: q<=8'b10100010;
	12'h0x105: q<=8'b10101010;
	12'h0x106: q<=8'b00100000;
	12'h0x107: q<=8'b01011010;
	12'h0x108: q<=8'b10110001;
	12'h0x109: q<=8'b10101101;
	12'h0x10a: q<=8'b01001110;
	12'h0x10b: q<=8'b00000001;
	12'h0x10c: q<=8'b11001001;
	12'h0x10d: q<=8'b10100000;
	12'h0x10e: q<=8'b10110000;
	12'h0x10f: q<=8'b00000101;
	12'h0x110: q<=8'b01101001;
	12'h0x111: q<=8'b00010100;
	12'h0x112: q<=8'b10001101;
	12'h0x113: q<=8'b01001110;
	12'h0x114: q<=8'b00000001;
	12'h0x115: q<=8'b11001001;
	12'h0x116: q<=8'b01010000;
	12'h0x117: q<=8'b10010000;
	12'h0x118: q<=8'b00010111;
	12'h0x119: q<=8'b10101101;
	12'h0x11a: q<=8'b01001101;
	12'h0x11b: q<=8'b00000001;
	12'h0x11c: q<=8'b00011000;
	12'h0x11d: q<=8'b01101001;
	12'h0x11e: q<=8'b00001000;
	12'h0x11f: q<=8'b10001101;
	12'h0x120: q<=8'b01001101;
	12'h0x121: q<=8'b00000001;
	12'h0x122: q<=8'b11001101;
	12'h0x123: q<=8'b01001110;
	12'h0x124: q<=8'b00000001;
	12'h0x125: q<=8'b10010000;
	12'h0x126: q<=8'b00001001;
	12'h0x127: q<=8'b10101001;
	12'h0x128: q<=8'b10100000;
	12'h0x129: q<=8'b10001101;
	12'h0x12a: q<=8'b01001101;
	12'h0x12b: q<=8'b00000001;
	12'h0x12c: q<=8'b10101001;
	12'h0x12d: q<=8'b00010100;
	12'h0x12e: q<=8'b10000101;
	12'h0x12f: q<=8'b00000001;
	12'h0x130: q<=8'b01100000;
	12'h0x131: q<=8'b10101001;
	12'h0x132: q<=8'b00111111;
	12'h0x133: q<=8'b10100010;
	12'h0x134: q<=8'b01001110;
	12'h0x135: q<=8'b00100000;
	12'h0x136: q<=8'b01011010;
	12'h0x137: q<=8'b10110001;
	12'h0x138: q<=8'b10101101;
	12'h0x139: q<=8'b01001101;
	12'h0x13a: q<=8'b00000001;
	12'h0x13b: q<=8'b11001001;
	12'h0x13c: q<=8'b00110000;
	12'h0x13d: q<=8'b10010000;
	12'h0x13e: q<=8'b00000101;
	12'h0x13f: q<=8'b11101001;
	12'h0x140: q<=8'b00000001;
	12'h0x141: q<=8'b10001101;
	12'h0x142: q<=8'b01001101;
	12'h0x143: q<=8'b00000001;
	12'h0x144: q<=8'b11001001;
	12'h0x145: q<=8'b10000000;
	12'h0x146: q<=8'b10110000;
	12'h0x147: q<=8'b00010001;
	12'h0x148: q<=8'b10101101;
	12'h0x149: q<=8'b01001110;
	12'h0x14a: q<=8'b00000001;
	12'h0x14b: q<=8'b00111000;
	12'h0x14c: q<=8'b11101001;
	12'h0x14d: q<=8'b00000001;
	12'h0x14e: q<=8'b11001101;
	12'h0x14f: q<=8'b01001101;
	12'h0x150: q<=8'b00000001;
	12'h0x151: q<=8'b10110000;
	12'h0x152: q<=8'b00000011;
	12'h0x153: q<=8'b10101101;
	12'h0x154: q<=8'b01001101;
	12'h0x155: q<=8'b00000001;
	12'h0x156: q<=8'b10001101;
	12'h0x157: q<=8'b01001110;
	12'h0x158: q<=8'b00000001;
	12'h0x159: q<=8'b01100000;
	12'h0x15a: q<=8'b10000101;
	12'h0x15b: q<=8'b01010111;
	12'h0x15c: q<=8'b10000110;
	12'h0x15d: q<=8'b01010110;
	12'h0x15e: q<=8'b10101101;
	12'h0x15f: q<=8'b01001101;
	12'h0x160: q<=8'b00000001;
	12'h0x161: q<=8'b10000101;
	12'h0x162: q<=8'b00110111;
	12'h0x163: q<=8'b11001110;
	12'h0x164: q<=8'b01101110;
	12'h0x165: q<=8'b00000001;
	12'h0x166: q<=8'b10100101;
	12'h0x167: q<=8'b00110111;
	12'h0x168: q<=8'b00001010;
	12'h0x169: q<=8'b00001010;
	12'h0x16a: q<=8'b00101001;
	12'h0x16b: q<=8'b01111111;
	12'h0x16c: q<=8'b10101000;
	12'h0x16d: q<=8'b10100101;
	12'h0x16e: q<=8'b00110111;
	12'h0x16f: q<=8'b01001010;
	12'h0x170: q<=8'b01001010;
	12'h0x171: q<=8'b01001010;
	12'h0x172: q<=8'b01001010;
	12'h0x173: q<=8'b01001010;
	12'h0x174: q<=8'b00100000;
	12'h0x175: q<=8'b01101100;
	12'h0x176: q<=8'b11011111;
	12'h0x177: q<=8'b10100101;
	12'h0x178: q<=8'b00110111;
	12'h0x179: q<=8'b11001101;
	12'h0x17a: q<=8'b01001101;
	12'h0x17b: q<=8'b00000001;
	12'h0x17c: q<=8'b11010000;
	12'h0x17d: q<=8'b00000101;
	12'h0x17e: q<=8'b10101001;
	12'h0x17f: q<=8'b00000000;
	12'h0x180: q<=8'b10111000;
	12'h0x181: q<=8'b01010000;
	12'h0x182: q<=8'b00001100;
	12'h0x183: q<=8'b01001010;
	12'h0x184: q<=8'b01001010;
	12'h0x185: q<=8'b01001010;
	12'h0x186: q<=8'b11101010;
	12'h0x187: q<=8'b00101001;
	12'h0x188: q<=8'b00000111;
	12'h0x189: q<=8'b11001001;
	12'h0x18a: q<=8'b00000111;
	12'h0x18b: q<=8'b11010000;
	12'h0x18c: q<=8'b00000010;
	12'h0x18d: q<=8'b10101001;
	12'h0x18e: q<=8'b00000011;
	12'h0x18f: q<=8'b10101000;
	12'h0x190: q<=8'b10101001;
	12'h0x191: q<=8'b01101000;
	12'h0x192: q<=8'b00100000;
	12'h0x193: q<=8'b01001100;
	12'h0x194: q<=8'b11011111;
	12'h0x195: q<=8'b10100101;
	12'h0x196: q<=8'b01010111;
	12'h0x197: q<=8'b10100110;
	12'h0x198: q<=8'b01010110;
	12'h0x199: q<=8'b00100000;
	12'h0x19a: q<=8'b00111001;
	12'h0x19b: q<=8'b11011111;
	12'h0x19c: q<=8'b10100101;
	12'h0x19d: q<=8'b00110111;
	12'h0x19e: q<=8'b00011000;
	12'h0x19f: q<=8'b01101001;
	12'h0x1a0: q<=8'b00000010;
	12'h0x1a1: q<=8'b10000101;
	12'h0x1a2: q<=8'b00110111;
	12'h0x1a3: q<=8'b11001101;
	12'h0x1a4: q<=8'b01001110;
	12'h0x1a5: q<=8'b00000001;
	12'h0x1a6: q<=8'b10010000;
	12'h0x1a7: q<=8'b10111110;
	12'h0x1a8: q<=8'b10100010;
	12'h0x1a9: q<=8'b00101100;
	12'h0x1aa: q<=8'b10101001;
	12'h0x1ab: q<=8'b11010000;
	12'h0x1ac: q<=8'b00100000;
	12'h0x1ad: q<=8'b00010111;
	12'h0x1ae: q<=8'b10101011;
	12'h0x1af: q<=8'b10101001;
	12'h0x1b0: q<=8'b00111111;
	12'h0x1b1: q<=8'b10100010;
	12'h0x1b2: q<=8'b11110010;
	12'h0x1b3: q<=8'b01001100;
	12'h0x1b4: q<=8'b00111001;
	12'h0x1b5: q<=8'b11011111;
	12'h0x1b6: q<=8'b00100000;
	12'h0x1b7: q<=8'b11000011;
	12'h0x1b8: q<=8'b11000001;
	12'h0x1b9: q<=8'b10101101;
	12'h0x1ba: q<=8'b00000000;
	12'h0x1bb: q<=8'b00100000;
	12'h0x1bc: q<=8'b11001101;
	12'h0x1bd: q<=8'b11000110;
	12'h0x1be: q<=8'b11001110;
	12'h0x1bf: q<=8'b11010000;
	12'h0x1c0: q<=8'b00000110;
	12'h0x1c1: q<=8'b10101101;
	12'h0x1c2: q<=8'b00110011;
	12'h0x1c3: q<=8'b00000001;
	12'h0x1c4: q<=8'b11010000;
	12'h0x1c5: q<=8'b00000001;
	12'h0x1c6: q<=8'b01100000;
	12'h0x1c7: q<=8'b10100101;
	12'h0x1c8: q<=8'b00000001;
	12'h0x1c9: q<=8'b11001001;
	12'h0x1ca: q<=8'b00000000;
	12'h0x1cb: q<=8'b11110000;
	12'h0x1cc: q<=8'b00111100;
	12'h0x1cd: q<=8'b10101001;
	12'h0x1ce: q<=8'b00000000;
	12'h0x1cf: q<=8'b00100000;
	12'h0x1d0: q<=8'b10111110;
	12'h0x1d1: q<=8'b10110010;
	12'h0x1d2: q<=8'b00100000;
	12'h0x1d3: q<=8'b00110010;
	12'h0x1d4: q<=8'b10110011;
	12'h0x1d5: q<=8'b10110000;
	12'h0x1d6: q<=8'b00011110;
	12'h0x1d7: q<=8'b00100000;
	12'h0x1d8: q<=8'b00001101;
	12'h0x1d9: q<=8'b10110010;
	12'h0x1da: q<=8'b10101101;
	12'h0x1db: q<=8'b01101110;
	12'h0x1dc: q<=8'b00000001;
	12'h0x1dd: q<=8'b11110000;
	12'h0x1de: q<=8'b00010110;
	12'h0x1df: q<=8'b10100000;
	12'h0x1e0: q<=8'b00100111;
	12'h0x1e1: q<=8'b10101001;
	12'h0x1e2: q<=8'b00001110;
	12'h0x1e3: q<=8'b00111000;
	12'h0x1e4: q<=8'b11110001;
	12'h0x1e5: q<=8'b10110110;
	12'h0x1e6: q<=8'b10001000;
	12'h0x1e7: q<=8'b00010000;
	12'h0x1e8: q<=8'b11111011;
	12'h0x1e9: q<=8'b10101000;
	12'h0x1ea: q<=8'b11110000;
	12'h0x1eb: q<=8'b00000010;
	12'h0x1ec: q<=8'b01001001;
	12'h0x1ed: q<=8'b11100101;
	12'h0x1ee: q<=8'b11110000;
	12'h0x1ef: q<=8'b00000010;
	12'h0x1f0: q<=8'b01001001;
	12'h0x1f1: q<=8'b00101001;
	12'h0x1f2: q<=8'b10001101;
	12'h0x1f3: q<=8'b01010101;
	12'h0x1f4: q<=8'b00000100;
	12'h0x1f5: q<=8'b10101001;
	12'h0x1f6: q<=8'b00000000;
	12'h0x1f7: q<=8'b00100000;
	12'h0x1f8: q<=8'b11111110;
	12'h0x1f9: q<=8'b10110010;
	12'h0x1fa: q<=8'b10101101;
	12'h0x1fb: q<=8'b11000100;
	12'h0x1fc: q<=8'b11001110;
	12'h0x1fd: q<=8'b10001101;
	12'h0x1fe: q<=8'b00000000;
	12'h0x1ff: q<=8'b00100000;
	12'h0x200: q<=8'b10101101;
	12'h0x201: q<=8'b11000101;
	12'h0x202: q<=8'b11001110;
	12'h0x203: q<=8'b10001101;
	12'h0x204: q<=8'b00000001;
	12'h0x205: q<=8'b00100000;
	12'h0x206: q<=8'b10111000;
	12'h0x207: q<=8'b01010000;
	12'h0x208: q<=8'b00000011;
	12'h0x209: q<=8'b01001100;
	12'h0x20a: q<=8'b00110000;
	12'h0x20b: q<=8'b10110010;
	12'h0x20c: q<=8'b01100000;
	12'h0x20d: q<=8'b10100110;
	12'h0x20e: q<=8'b00000001;
	12'h0x20f: q<=8'b10111101;
	12'h0x210: q<=8'b00011001;
	12'h0x211: q<=8'b10110010;
	12'h0x212: q<=8'b01001000;
	12'h0x213: q<=8'b10111101;
	12'h0x214: q<=8'b00011000;
	12'h0x215: q<=8'b10110010;
	12'h0x216: q<=8'b01001000;
	12'h0x217: q<=8'b01100000;
	12'h0x218: q<=8'b00101111;
	12'h0x219: q<=8'b10110010;
	12'h0x21a: q<=8'b00000011;
	12'h0x21b: q<=8'b11011000;
	12'h0x21c: q<=8'b10111001;
	12'h0x21d: q<=8'b10111000;
	12'h0x21e: q<=8'b11101001;
	12'h0x21f: q<=8'b10101101;
	12'h0x220: q<=8'b10000000;
	12'h0x221: q<=8'b10101111;
	12'h0x222: q<=8'b00011011;
	12'h0x223: q<=8'b10101110;
	12'h0x224: q<=8'b01100001;
	12'h0x225: q<=8'b10101010;
	12'h0x226: q<=8'b01011001;
	12'h0x227: q<=8'b10101010;
	12'h0x228: q<=8'b01101110;
	12'h0x229: q<=8'b10101010;
	12'h0x22a: q<=8'b00000001;
	12'h0x22b: q<=8'b10110001;
	12'h0x22c: q<=8'b00110000;
	12'h0x22d: q<=8'b10110001;
	12'h0x22e: q<=8'b01111000;
	12'h0x22f: q<=8'b10101010;
	12'h0x230: q<=8'b10101001;
	12'h0x231: q<=8'b00000111;
	12'h0x232: q<=8'b00100000;
	12'h0x233: q<=8'b10111110;
	12'h0x234: q<=8'b10110010;
	12'h0x235: q<=8'b00100000;
	12'h0x236: q<=8'b10000110;
	12'h0x237: q<=8'b10110101;
	12'h0x238: q<=8'b10101001;
	12'h0x239: q<=8'b00000111;
	12'h0x23a: q<=8'b00100000;
	12'h0x23b: q<=8'b11111110;
	12'h0x23c: q<=8'b10110010;
	12'h0x23d: q<=8'b10101001;
	12'h0x23e: q<=8'b00000100;
	12'h0x23f: q<=8'b00100000;
	12'h0x240: q<=8'b10111110;
	12'h0x241: q<=8'b10110010;
	12'h0x242: q<=8'b00100000;
	12'h0x243: q<=8'b01011011;
	12'h0x244: q<=8'b10110111;
	12'h0x245: q<=8'b10101001;
	12'h0x246: q<=8'b00000100;
	12'h0x247: q<=8'b00100000;
	12'h0x248: q<=8'b11111110;
	12'h0x249: q<=8'b10110010;
	12'h0x24a: q<=8'b10101001;
	12'h0x24b: q<=8'b00000011;
	12'h0x24c: q<=8'b00100000;
	12'h0x24d: q<=8'b10111110;
	12'h0x24e: q<=8'b10110010;
	12'h0x24f: q<=8'b00100000;
	12'h0x250: q<=8'b10101101;
	12'h0x251: q<=8'b10110101;
	12'h0x252: q<=8'b10101001;
	12'h0x253: q<=8'b00000011;
	12'h0x254: q<=8'b00100000;
	12'h0x255: q<=8'b11111110;
	12'h0x256: q<=8'b10110010;
	12'h0x257: q<=8'b10101001;
	12'h0x258: q<=8'b00000110;
	12'h0x259: q<=8'b00100000;
	12'h0x25a: q<=8'b10111110;
	12'h0x25b: q<=8'b10110010;
	12'h0x25c: q<=8'b00100000;
	12'h0x25d: q<=8'b10011010;
	12'h0x25e: q<=8'b10110111;
	12'h0x25f: q<=8'b10101001;
	12'h0x260: q<=8'b00000110;
	12'h0x261: q<=8'b00100000;
	12'h0x262: q<=8'b11111110;
	12'h0x263: q<=8'b10110010;
	12'h0x264: q<=8'b10101001;
	12'h0x265: q<=8'b00000101;
	12'h0x266: q<=8'b00100000;
	12'h0x267: q<=8'b10111110;
	12'h0x268: q<=8'b10110010;
	12'h0x269: q<=8'b00100000;
	12'h0x26a: q<=8'b10011000;
	12'h0x26b: q<=8'b10110100;
	12'h0x26c: q<=8'b10101001;
	12'h0x26d: q<=8'b00000101;
	12'h0x26e: q<=8'b00100000;
	12'h0x26f: q<=8'b11111110;
	12'h0x270: q<=8'b10110010;
	12'h0x271: q<=8'b10101001;
	12'h0x272: q<=8'b00000000;
	12'h0x273: q<=8'b00100000;
	12'h0x274: q<=8'b10111110;
	12'h0x275: q<=8'b10110010;
	12'h0x276: q<=8'b00100000;
	12'h0x277: q<=8'b10110100;
	12'h0x278: q<=8'b10101000;
	12'h0x279: q<=8'b10100101;
	12'h0x27a: q<=8'b00000101;
	12'h0x27b: q<=8'b00110000;
	12'h0x27c: q<=8'b00001101;
	12'h0x27d: q<=8'b10101001;
	12'h0x27e: q<=8'b11110010;
	12'h0x27f: q<=8'b00011000;
	12'h0x280: q<=8'b10100000;
	12'h0x281: q<=8'b00100111;
	12'h0x282: q<=8'b01110001;
	12'h0x283: q<=8'b10110110;
	12'h0x284: q<=8'b10001000;
	12'h0x285: q<=8'b00010000;
	12'h0x286: q<=8'b11111011;
	12'h0x287: q<=8'b10001101;
	12'h0x288: q<=8'b00011011;
	12'h0x289: q<=8'b00000001;
	12'h0x28a: q<=8'b10101001;
	12'h0x28b: q<=8'b00000000;
	12'h0x28c: q<=8'b00100000;
	12'h0x28d: q<=8'b11111110;
	12'h0x28e: q<=8'b10110010;
	12'h0x28f: q<=8'b00100000;
	12'h0x290: q<=8'b01100111;
	12'h0x291: q<=8'b10110011;
	12'h0x292: q<=8'b10101001;
	12'h0x293: q<=8'b00000001;
	12'h0x294: q<=8'b00100000;
	12'h0x295: q<=8'b10111110;
	12'h0x296: q<=8'b10110010;
	12'h0x297: q<=8'b00100000;
	12'h0x298: q<=8'b11000010;
	12'h0x299: q<=8'b11000101;
	12'h0x29a: q<=8'b10101001;
	12'h0x29b: q<=8'b00000001;
	12'h0x29c: q<=8'b00100000;
	12'h0x29d: q<=8'b11111110;
	12'h0x29e: q<=8'b10110010;
	12'h0x29f: q<=8'b10101001;
	12'h0x2a0: q<=8'b00001000;
	12'h0x2a1: q<=8'b00100000;
	12'h0x2a2: q<=8'b10111110;
	12'h0x2a3: q<=8'b10110010;
	12'h0x2a4: q<=8'b00100000;
	12'h0x2a5: q<=8'b01001101;
	12'h0x2a6: q<=8'b11000101;
	12'h0x2a7: q<=8'b10101001;
	12'h0x2a8: q<=8'b00001000;
	12'h0x2a9: q<=8'b00100000;
	12'h0x2aa: q<=8'b11111110;
	12'h0x2ab: q<=8'b10110010;
	12'h0x2ac: q<=8'b10101001;
	12'h0x2ad: q<=8'b00000000;
	12'h0x2ae: q<=8'b10001101;
	12'h0x2af: q<=8'b00010100;
	12'h0x2b0: q<=8'b00000001;
	12'h0x2b1: q<=8'b10101101;
	12'h0x2b2: q<=8'b11000010;
	12'h0x2b3: q<=8'b11001110;
	12'h0x2b4: q<=8'b10001101;
	12'h0x2b5: q<=8'b00000000;
	12'h0x2b6: q<=8'b00100000;
	12'h0x2b7: q<=8'b10101101;
	12'h0x2b8: q<=8'b11000011;
	12'h0x2b9: q<=8'b11001110;
	12'h0x2ba: q<=8'b10001101;
	12'h0x2bb: q<=8'b00000001;
	12'h0x2bc: q<=8'b00100000;
	12'h0x2bd: q<=8'b01100000;
	12'h0x2be: q<=8'b10101010;
	12'h0x2bf: q<=8'b00001010;
	12'h0x2c0: q<=8'b10101000;
	12'h0x2c1: q<=8'b10111101;
	12'h0x2c2: q<=8'b00010101;
	12'h0x2c3: q<=8'b00000100;
	12'h0x2c4: q<=8'b11010000;
	12'h0x2c5: q<=8'b00001001;
	12'h0x2c6: q<=8'b10111110;
	12'h0x2c7: q<=8'b01111010;
	12'h0x2c8: q<=8'b11001110;
	12'h0x2c9: q<=8'b10111001;
	12'h0x2ca: q<=8'b01111011;
	12'h0x2cb: q<=8'b11001110;
	12'h0x2cc: q<=8'b10111000;
	12'h0x2cd: q<=8'b01010000;
	12'h0x2ce: q<=8'b00000110;
	12'h0x2cf: q<=8'b10111110;
	12'h0x2d0: q<=8'b01101000;
	12'h0x2d1: q<=8'b11001110;
	12'h0x2d2: q<=8'b10111001;
	12'h0x2d3: q<=8'b01101001;
	12'h0x2d4: q<=8'b11001110;
	12'h0x2d5: q<=8'b10000110;
	12'h0x2d6: q<=8'b01110100;
	12'h0x2d7: q<=8'b10000101;
	12'h0x2d8: q<=8'b01110101;
	12'h0x2d9: q<=8'b10101001;
	12'h0x2da: q<=8'b00000000;
	12'h0x2db: q<=8'b10000101;
	12'h0x2dc: q<=8'b10101001;
	12'h0x2dd: q<=8'b01100000;
	12'h0x2de: q<=8'b10101010;
	12'h0x2df: q<=8'b00001010;
	12'h0x2e0: q<=8'b10101000;
	12'h0x2e1: q<=8'b10111101;
	12'h0x2e2: q<=8'b00010101;
	12'h0x2e3: q<=8'b00000100;
	12'h0x2e4: q<=8'b11010000;
	12'h0x2e5: q<=8'b00001001;
	12'h0x2e6: q<=8'b10111110;
	12'h0x2e7: q<=8'b01101000;
	12'h0x2e8: q<=8'b11001110;
	12'h0x2e9: q<=8'b10111001;
	12'h0x2ea: q<=8'b01101001;
	12'h0x2eb: q<=8'b11001110;
	12'h0x2ec: q<=8'b10111000;
	12'h0x2ed: q<=8'b01010000;
	12'h0x2ee: q<=8'b00000110;
	12'h0x2ef: q<=8'b10111110;
	12'h0x2f0: q<=8'b01111010;
	12'h0x2f1: q<=8'b11001110;
	12'h0x2f2: q<=8'b10111001;
	12'h0x2f3: q<=8'b01111011;
	12'h0x2f4: q<=8'b11001110;
	12'h0x2f5: q<=8'b10000110;
	12'h0x2f6: q<=8'b00111011;
	12'h0x2f7: q<=8'b10000101;
	12'h0x2f8: q<=8'b00111100;
	12'h0x2f9: q<=8'b10101001;
	12'h0x2fa: q<=8'b00000000;
	12'h0x2fb: q<=8'b10000101;
	12'h0x2fc: q<=8'b10101001;
	12'h0x2fd: q<=8'b01100000;
	12'h0x2fe: q<=8'b01001000;
	12'h0x2ff: q<=8'b00100000;
	12'h0x300: q<=8'b00001001;
	12'h0x301: q<=8'b11011111;
	12'h0x302: q<=8'b01101000;
	12'h0x303: q<=8'b10101010;
	12'h0x304: q<=8'b00001010;
	12'h0x305: q<=8'b10101000;
	12'h0x306: q<=8'b10111001;
	12'h0x307: q<=8'b10001100;
	12'h0x308: q<=8'b11001110;
	12'h0x309: q<=8'b10000101;
	12'h0x30a: q<=8'b00111011;
	12'h0x30b: q<=8'b10111001;
	12'h0x30c: q<=8'b10001101;
	12'h0x30d: q<=8'b11001110;
	12'h0x30e: q<=8'b10000101;
	12'h0x30f: q<=8'b00111100;
	12'h0x310: q<=8'b10111101;
	12'h0x311: q<=8'b00010101;
	12'h0x312: q<=8'b00000100;
	12'h0x313: q<=8'b01001001;
	12'h0x314: q<=8'b00000001;
	12'h0x315: q<=8'b10011101;
	12'h0x316: q<=8'b00010101;
	12'h0x317: q<=8'b00000100;
	12'h0x318: q<=8'b11010000;
	12'h0x319: q<=8'b00001001;
	12'h0x31a: q<=8'b10111001;
	12'h0x31b: q<=8'b10011110;
	12'h0x31c: q<=8'b11001110;
	12'h0x31d: q<=8'b10111110;
	12'h0x31e: q<=8'b10011111;
	12'h0x31f: q<=8'b11001110;
	12'h0x320: q<=8'b10111000;
	12'h0x321: q<=8'b01010000;
	12'h0x322: q<=8'b00000110;
	12'h0x323: q<=8'b10111001;
	12'h0x324: q<=8'b10110000;
	12'h0x325: q<=8'b11001110;
	12'h0x326: q<=8'b10111110;
	12'h0x327: q<=8'b10110001;
	12'h0x328: q<=8'b11001110;
	12'h0x329: q<=8'b10100000;
	12'h0x32a: q<=8'b00000000;
	12'h0x32b: q<=8'b10010001;
	12'h0x32c: q<=8'b00111011;
	12'h0x32d: q<=8'b10001010;
	12'h0x32e: q<=8'b11001000;
	12'h0x32f: q<=8'b10010001;
	12'h0x330: q<=8'b00111011;
	12'h0x331: q<=8'b01100000;
	12'h0x332: q<=8'b10101101;
	12'h0x333: q<=8'b11000100;
	12'h0x334: q<=8'b11001110;
	12'h0x335: q<=8'b11001101;
	12'h0x336: q<=8'b00000000;
	12'h0x337: q<=8'b00100000;
	12'h0x338: q<=8'b11110000;
	12'h0x339: q<=8'b00000101;
	12'h0x33a: q<=8'b10001101;
	12'h0x33b: q<=8'b00000000;
	12'h0x33c: q<=8'b00100000;
	12'h0x33d: q<=8'b00111000;
	12'h0x33e: q<=8'b01100000;
	12'h0x33f: q<=8'b10101101;
	12'h0x340: q<=8'b00010101;
	12'h0x341: q<=8'b00000100;
	12'h0x342: q<=8'b11010000;
	12'h0x343: q<=8'b00000101;
	12'h0x344: q<=8'b10100010;
	12'h0x345: q<=8'b00000010;
	12'h0x346: q<=8'b10111000;
	12'h0x347: q<=8'b01010000;
	12'h0x348: q<=8'b00000010;
	12'h0x349: q<=8'b10100010;
	12'h0x34a: q<=8'b00001000;
	12'h0x34b: q<=8'b10111101;
	12'h0x34c: q<=8'b10011110;
	12'h0x34d: q<=8'b11001110;
	12'h0x34e: q<=8'b10100000;
	12'h0x34f: q<=8'b00000000;
	12'h0x350: q<=8'b10001100;
	12'h0x351: q<=8'b01101110;
	12'h0x352: q<=8'b00000001;
	12'h0x353: q<=8'b10010001;
	12'h0x354: q<=8'b01110100;
	12'h0x355: q<=8'b11001000;
	12'h0x356: q<=8'b10111101;
	12'h0x357: q<=8'b10011111;
	12'h0x358: q<=8'b11001110;
	12'h0x359: q<=8'b10010001;
	12'h0x35a: q<=8'b01110100;
	12'h0x35b: q<=8'b10111101;
	12'h0x35c: q<=8'b01101000;
	12'h0x35d: q<=8'b11001110;
	12'h0x35e: q<=8'b10000101;
	12'h0x35f: q<=8'b01110100;
	12'h0x360: q<=8'b10111101;
	12'h0x361: q<=8'b01101001;
	12'h0x362: q<=8'b11001110;
	12'h0x363: q<=8'b10000101;
	12'h0x364: q<=8'b01110101;
	12'h0x365: q<=8'b00011000;
	12'h0x366: q<=8'b01100000;
	12'h0x367: q<=8'b10101101;
	12'h0x368: q<=8'b00010100;
	12'h0x369: q<=8'b00000001;
	12'h0x36a: q<=8'b11110000;
	12'h0x36b: q<=8'b00001101;
	12'h0x36c: q<=8'b10101001;
	12'h0x36d: q<=8'b00000010;
	12'h0x36e: q<=8'b00100000;
	12'h0x36f: q<=8'b10111110;
	12'h0x370: q<=8'b10110010;
	12'h0x371: q<=8'b00100000;
	12'h0x372: q<=8'b00001101;
	12'h0x373: q<=8'b11000011;
	12'h0x374: q<=8'b10101001;
	12'h0x375: q<=8'b00000010;
	12'h0x376: q<=8'b00100000;
	12'h0x377: q<=8'b11111110;
	12'h0x378: q<=8'b10110010;
	12'h0x379: q<=8'b10101001;
	12'h0x37a: q<=8'b00000010;
	12'h0x37b: q<=8'b00100000;
	12'h0x37c: q<=8'b11011110;
	12'h0x37d: q<=8'b10110010;
	12'h0x37e: q<=8'b10101001;
	12'h0x37f: q<=8'b00000000;
	12'h0x380: q<=8'b10100010;
	12'h0x381: q<=8'b00001111;
	12'h0x382: q<=8'b10011101;
	12'h0x383: q<=8'b00100101;
	12'h0x384: q<=8'b00000100;
	12'h0x385: q<=8'b11001010;
	12'h0x386: q<=8'b00010000;
	12'h0x387: q<=8'b11111010;
	12'h0x388: q<=8'b10101101;
	12'h0x389: q<=8'b00000110;
	12'h0x38a: q<=8'b00000001;
	12'h0x38b: q<=8'b00110000;
	12'h0x38c: q<=8'b01001001;
	12'h0x38d: q<=8'b10101110;
	12'h0x38e: q<=8'b00011100;
	12'h0x38f: q<=8'b00000001;
	12'h0x390: q<=8'b10111101;
	12'h0x391: q<=8'b11011111;
	12'h0x392: q<=8'b00000010;
	12'h0x393: q<=8'b11110000;
	12'h0x394: q<=8'b00111110;
	12'h0x395: q<=8'b10100000;
	12'h0x396: q<=8'b00000000;
	12'h0x397: q<=8'b10111101;
	12'h0x398: q<=8'b10000011;
	12'h0x399: q<=8'b00000010;
	12'h0x39a: q<=8'b00101001;
	12'h0x39b: q<=8'b00000111;
	12'h0x39c: q<=8'b11001001;
	12'h0x39d: q<=8'b00000001;
	12'h0x39e: q<=8'b11010000;
	12'h0x39f: q<=8'b00110011;
	12'h0x3a0: q<=8'b11001000;
	12'h0x3a1: q<=8'b10000100;
	12'h0x3a2: q<=8'b00101001;
	12'h0x3a3: q<=8'b10111101;
	12'h0x3a4: q<=8'b10000011;
	12'h0x3a5: q<=8'b00000010;
	12'h0x3a6: q<=8'b00101001;
	12'h0x3a7: q<=8'b10000000;
	12'h0x3a8: q<=8'b11010000;
	12'h0x3a9: q<=8'b00011100;
	12'h0x3aa: q<=8'b10101101;
	12'h0x3ab: q<=8'b01001000;
	12'h0x3ac: q<=8'b00000001;
	12'h0x3ad: q<=8'b00110000;
	12'h0x3ae: q<=8'b00001100;
	12'h0x3af: q<=8'b10111101;
	12'h0x3b0: q<=8'b11011111;
	12'h0x3b1: q<=8'b00000010;
	12'h0x3b2: q<=8'b11001101;
	12'h0x3b3: q<=8'b01010111;
	12'h0x3b4: q<=8'b00000001;
	12'h0x3b5: q<=8'b10110000;
	12'h0x3b6: q<=8'b00000100;
	12'h0x3b7: q<=8'b11100110;
	12'h0x3b8: q<=8'b00101001;
	12'h0x3b9: q<=8'b11100110;
	12'h0x3ba: q<=8'b00101001;
	12'h0x3bb: q<=8'b10100101;
	12'h0x3bc: q<=8'b00101001;
	12'h0x3bd: q<=8'b10111100;
	12'h0x3be: q<=8'b11001100;
	12'h0x3bf: q<=8'b00000010;
	12'h0x3c0: q<=8'b00011001;
	12'h0x3c1: q<=8'b00100101;
	12'h0x3c2: q<=8'b00000100;
	12'h0x3c3: q<=8'b10011001;
	12'h0x3c4: q<=8'b00100101;
	12'h0x3c5: q<=8'b00000100;
	12'h0x3c6: q<=8'b10111100;
	12'h0x3c7: q<=8'b10111001;
	12'h0x3c8: q<=8'b00000010;
	12'h0x3c9: q<=8'b10100101;
	12'h0x3ca: q<=8'b00101001;
	12'h0x3cb: q<=8'b00001001;
	12'h0x3cc: q<=8'b10000000;
	12'h0x3cd: q<=8'b00011001;
	12'h0x3ce: q<=8'b00100101;
	12'h0x3cf: q<=8'b00000100;
	12'h0x3d0: q<=8'b10011001;
	12'h0x3d1: q<=8'b00100101;
	12'h0x3d2: q<=8'b00000100;
	12'h0x3d3: q<=8'b11001010;
	12'h0x3d4: q<=8'b00010000;
	12'h0x3d5: q<=8'b10111010;
	12'h0x3d6: q<=8'b10101001;
	12'h0x3d7: q<=8'b00000110;
	12'h0x3d8: q<=8'b10101100;
	12'h0x3d9: q<=8'b00100101;
	12'h0x3da: q<=8'b00000001;
	12'h0x3db: q<=8'b11110000;
	12'h0x3dc: q<=8'b00001100;
	12'h0x3dd: q<=8'b00110000;
	12'h0x3de: q<=8'b00001010;
	12'h0x3df: q<=8'b10100101;
	12'h0x3e0: q<=8'b00000011;
	12'h0x3e1: q<=8'b00101001;
	12'h0x3e2: q<=8'b00000111;
	12'h0x3e3: q<=8'b11001001;
	12'h0x3e4: q<=8'b00000111;
	12'h0x3e5: q<=8'b11010000;
	12'h0x3e6: q<=8'b00000010;
	12'h0x3e7: q<=8'b10101001;
	12'h0x3e8: q<=8'b00000001;
	12'h0x3e9: q<=8'b10000101;
	12'h0x3ea: q<=8'b00101001;
	12'h0x3eb: q<=8'b10100000;
	12'h0x3ec: q<=8'b11111111;
	12'h0x3ed: q<=8'b10100010;
	12'h0x3ee: q<=8'b11111111;
	12'h0x3ef: q<=8'b10000110;
	12'h0x3f0: q<=8'b00101100;
	12'h0x3f1: q<=8'b10101101;
	12'h0x3f2: q<=8'b00000010;
	12'h0x3f3: q<=8'b00000010;
	12'h0x3f4: q<=8'b11110000;
	12'h0x3f5: q<=8'b00001011;
	12'h0x3f6: q<=8'b10101101;
	12'h0x3f7: q<=8'b00000001;
	12'h0x3f8: q<=8'b00000010;
	12'h0x3f9: q<=8'b00110000;
	12'h0x3fa: q<=8'b00000110;
	12'h0x3fb: q<=8'b10101110;
	12'h0x3fc: q<=8'b00000000;
	12'h0x3fd: q<=8'b00000010;
	12'h0x3fe: q<=8'b10101100;
	12'h0x3ff: q<=8'b00000001;
	12'h0x400: q<=8'b00000010;
	12'h0x401: q<=8'b10000110;
	12'h0x402: q<=8'b00101010;
	12'h0x403: q<=8'b10000100;
	12'h0x404: q<=8'b00101011;
	12'h0x405: q<=8'b10101101;
	12'h0x406: q<=8'b00100100;
	12'h0x407: q<=8'b00000001;
	12'h0x408: q<=8'b00110000;
	12'h0x409: q<=8'b00001000;
	12'h0x40a: q<=8'b00101001;
	12'h0x40b: q<=8'b00001110;
	12'h0x40c: q<=8'b01001010;
	12'h0x40d: q<=8'b10000101;
	12'h0x40e: q<=8'b00101100;
	12'h0x40f: q<=8'b11001110;
	12'h0x410: q<=8'b00100100;
	12'h0x411: q<=8'b00000001;
	12'h0x412: q<=8'b10100010;
	12'h0x413: q<=8'b00001111;
	12'h0x414: q<=8'b10100000;
	12'h0x415: q<=8'b00000110;
	12'h0x416: q<=8'b10111101;
	12'h0x417: q<=8'b00100101;
	12'h0x418: q<=8'b00000100;
	12'h0x419: q<=8'b11110000;
	12'h0x41a: q<=8'b00001100;
	12'h0x41b: q<=8'b00101001;
	12'h0x41c: q<=8'b00000010;
	12'h0x41d: q<=8'b11110000;
	12'h0x41e: q<=8'b00000101;
	12'h0x41f: q<=8'b10100101;
	12'h0x420: q<=8'b00000011;
	12'h0x421: q<=8'b00101001;
	12'h0x422: q<=8'b00000001;
	12'h0x423: q<=8'b10101000;
	12'h0x424: q<=8'b10111000;
	12'h0x425: q<=8'b01010000;
	12'h0x426: q<=8'b00100100;
	12'h0x427: q<=8'b11100100;
	12'h0x428: q<=8'b00101010;
	12'h0x429: q<=8'b11110000;
	12'h0x42a: q<=8'b00000010;
	12'h0x42b: q<=8'b11100100;
	12'h0x42c: q<=8'b00101011;
	12'h0x42d: q<=8'b11010000;
	12'h0x42e: q<=8'b00000101;
	12'h0x42f: q<=8'b10100000;
	12'h0x430: q<=8'b00000001;
	12'h0x431: q<=8'b10111000;
	12'h0x432: q<=8'b01010000;
	12'h0x433: q<=8'b00010111;
	12'h0x434: q<=8'b10101101;
	12'h0x435: q<=8'b00100100;
	12'h0x436: q<=8'b00000001;
	12'h0x437: q<=8'b00110000;
	12'h0x438: q<=8'b00010000;
	12'h0x439: q<=8'b10001010;
	12'h0x43a: q<=8'b00011000;
	12'h0x43b: q<=8'b01100101;
	12'h0x43c: q<=8'b00101100;
	12'h0x43d: q<=8'b00101001;
	12'h0x43e: q<=8'b00000111;
	12'h0x43f: q<=8'b11001001;
	12'h0x440: q<=8'b00000111;
	12'h0x441: q<=8'b11010000;
	12'h0x442: q<=8'b00000010;
	12'h0x443: q<=8'b10101001;
	12'h0x444: q<=8'b00000011;
	12'h0x445: q<=8'b10101000;
	12'h0x446: q<=8'b10111000;
	12'h0x447: q<=8'b01010000;
	12'h0x448: q<=8'b00000010;
	12'h0x449: q<=8'b10100100;
	12'h0x44a: q<=8'b00101001;
	12'h0x44b: q<=8'b10011000;
	12'h0x44c: q<=8'b10111100;
	12'h0x44d: q<=8'b01110110;
	12'h0x44e: q<=8'b10110100;
	12'h0x44f: q<=8'b10010001;
	12'h0x450: q<=8'b00111011;
	12'h0x451: q<=8'b11001010;
	12'h0x452: q<=8'b00010000;
	12'h0x453: q<=8'b11000000;
	12'h0x454: q<=8'b10100010;
	12'h0x455: q<=8'b00001111;
	12'h0x456: q<=8'b00101100;
	12'h0x457: q<=8'b00010001;
	12'h0x458: q<=8'b00000001;
	12'h0x459: q<=8'b00010000;
	12'h0x45a: q<=8'b00000001;
	12'h0x45b: q<=8'b11001010;
	12'h0x45c: q<=8'b10100000;
	12'h0x45d: q<=8'b11000000;
	12'h0x45e: q<=8'b10111101;
	12'h0x45f: q<=8'b00100101;
	12'h0x460: q<=8'b00000100;
	12'h0x461: q<=8'b00010000;
	12'h0x462: q<=8'b00000010;
	12'h0x463: q<=8'b10100000;
	12'h0x464: q<=8'b00000000;
	12'h0x465: q<=8'b10000100;
	12'h0x466: q<=8'b01011000;
	12'h0x467: q<=8'b10111100;
	12'h0x468: q<=8'b10000111;
	12'h0x469: q<=8'b10110100;
	12'h0x46a: q<=8'b10110001;
	12'h0x46b: q<=8'b10110000;
	12'h0x46c: q<=8'b00101001;
	12'h0x46d: q<=8'b00011111;
	12'h0x46e: q<=8'b00000101;
	12'h0x46f: q<=8'b01011000;
	12'h0x470: q<=8'b10010001;
	12'h0x471: q<=8'b10110000;
	12'h0x472: q<=8'b11001010;
	12'h0x473: q<=8'b00010000;
	12'h0x474: q<=8'b11100111;
	12'h0x475: q<=8'b01100000;
	12'h0x476: q<=8'b10101000;
	12'h0x477: q<=8'b10011100;
	12'h0x478: q<=8'b10010010;
	12'h0x479: q<=8'b10000110;
	12'h0x47a: q<=8'b01111100;
	12'h0x47b: q<=8'b01110000;
	12'h0x47c: q<=8'b01100110;
	12'h0x47d: q<=8'b01011010;
	12'h0x47e: q<=8'b01010000;
	12'h0x47f: q<=8'b01000100;
	12'h0x480: q<=8'b00111010;
	12'h0x481: q<=8'b00101110;
	12'h0x482: q<=8'b00100100;
	12'h0x483: q<=8'b00011000;
	12'h0x484: q<=8'b00001110;
	12'h0x485: q<=8'b00000010;
	12'h0x486: q<=8'b10110010;
	12'h0x487: q<=8'b00111011;
	12'h0x488: q<=8'b00110111;
	12'h0x489: q<=8'b00110011;
	12'h0x48a: q<=8'b00101111;
	12'h0x48b: q<=8'b00101011;
	12'h0x48c: q<=8'b00100111;
	12'h0x48d: q<=8'b00100011;
	12'h0x48e: q<=8'b00011111;
	12'h0x48f: q<=8'b00011011;
	12'h0x490: q<=8'b00010111;
	12'h0x491: q<=8'b00010011;
	12'h0x492: q<=8'b00001111;
	12'h0x493: q<=8'b00001011;
	12'h0x494: q<=8'b00000111;
	12'h0x495: q<=8'b00000011;
	12'h0x496: q<=8'b00111111;
	12'h0x497: q<=8'b00011101;
	12'h0x498: q<=8'b10100000;
	12'h0x499: q<=8'b00001100;
	12'h0x49a: q<=8'b10000100;
	12'h0x49b: q<=8'b10011110;
	12'h0x49c: q<=8'b10101001;
	12'h0x49d: q<=8'b00001000;
	12'h0x49e: q<=8'b00100000;
	12'h0x49f: q<=8'b01001100;
	12'h0x4a0: q<=8'b11011111;
	12'h0x4a1: q<=8'b10100010;
	12'h0x4a2: q<=8'b01100110;
	12'h0x4a3: q<=8'b00100000;
	12'h0x4a4: q<=8'b01100101;
	12'h0x4a5: q<=8'b11000111;
	12'h0x4a6: q<=8'b10101001;
	12'h0x4a7: q<=8'b00010010;
	12'h0x4a8: q<=8'b10000101;
	12'h0x4a9: q<=8'b01010110;
	12'h0x4aa: q<=8'b10100010;
	12'h0x4ab: q<=8'b00111111;
	12'h0x4ac: q<=8'b10000110;
	12'h0x4ad: q<=8'b00110111;
	12'h0x4ae: q<=8'b10100000;
	12'h0x4af: q<=8'b00000000;
	12'h0x4b0: q<=8'b10100110;
	12'h0x4b1: q<=8'b00110111;
	12'h0x4b2: q<=8'b10111101;
	12'h0x4b3: q<=8'b01000011;
	12'h0x4b4: q<=8'b00000010;
	12'h0x4b5: q<=8'b11010000;
	12'h0x4b6: q<=8'b00000011;
	12'h0x4b7: q<=8'b01001100;
	12'h0x4b8: q<=8'b01001001;
	12'h0x4b9: q<=8'b10110101;
	12'h0x4ba: q<=8'b11001001;
	12'h0x4bb: q<=8'b01010000;
	12'h0x4bc: q<=8'b10010000;
	12'h0x4bd: q<=8'b00000010;
	12'h0x4be: q<=8'b11000110;
	12'h0x4bf: q<=8'b00110111;
	12'h0x4c0: q<=8'b01001000;
	12'h0x4c1: q<=8'b00101001;
	12'h0x4c2: q<=8'b00111111;
	12'h0x4c3: q<=8'b10010001;
	12'h0x4c4: q<=8'b01110100;
	12'h0x4c5: q<=8'b01101000;
	12'h0x4c6: q<=8'b00101010;
	12'h0x4c7: q<=8'b00101010;
	12'h0x4c8: q<=8'b00101010;
	12'h0x4c9: q<=8'b00101001;
	12'h0x4ca: q<=8'b00000011;
	12'h0x4cb: q<=8'b00011000;
	12'h0x4cc: q<=8'b01101001;
	12'h0x4cd: q<=8'b00000001;
	12'h0x4ce: q<=8'b00001001;
	12'h0x4cf: q<=8'b01110000;
	12'h0x4d0: q<=8'b11001000;
	12'h0x4d1: q<=8'b10010001;
	12'h0x4d2: q<=8'b01110100;
	12'h0x4d3: q<=8'b11001000;
	12'h0x4d4: q<=8'b10111101;
	12'h0x4d5: q<=8'b00000011;
	12'h0x4d6: q<=8'b00000010;
	12'h0x4d7: q<=8'b10101010;
	12'h0x4d8: q<=8'b10111101;
	12'h0x4d9: q<=8'b10001010;
	12'h0x4da: q<=8'b00000011;
	12'h0x4db: q<=8'b00111000;
	12'h0x4dc: q<=8'b11100101;
	12'h0x4dd: q<=8'b01101000;
	12'h0x4de: q<=8'b10000101;
	12'h0x4df: q<=8'b01100011;
	12'h0x4e0: q<=8'b10010001;
	12'h0x4e1: q<=8'b01110100;
	12'h0x4e2: q<=8'b11001000;
	12'h0x4e3: q<=8'b10111101;
	12'h0x4e4: q<=8'b01111010;
	12'h0x4e5: q<=8'b00000011;
	12'h0x4e6: q<=8'b11100101;
	12'h0x4e7: q<=8'b01101001;
	12'h0x4e8: q<=8'b10000101;
	12'h0x4e9: q<=8'b01100100;
	12'h0x4ea: q<=8'b00101001;
	12'h0x4eb: q<=8'b00011111;
	12'h0x4ec: q<=8'b10010001;
	12'h0x4ed: q<=8'b01110100;
	12'h0x4ee: q<=8'b11001000;
	12'h0x4ef: q<=8'b10111101;
	12'h0x4f0: q<=8'b01101010;
	12'h0x4f1: q<=8'b00000011;
	12'h0x4f2: q<=8'b10000101;
	12'h0x4f3: q<=8'b01100001;
	12'h0x4f4: q<=8'b10010001;
	12'h0x4f5: q<=8'b01110100;
	12'h0x4f6: q<=8'b11001000;
	12'h0x4f7: q<=8'b10111101;
	12'h0x4f8: q<=8'b01011010;
	12'h0x4f9: q<=8'b00000011;
	12'h0x4fa: q<=8'b10000101;
	12'h0x4fb: q<=8'b01100010;
	12'h0x4fc: q<=8'b00101001;
	12'h0x4fd: q<=8'b00011111;
	12'h0x4fe: q<=8'b10010001;
	12'h0x4ff: q<=8'b01110100;
	12'h0x500: q<=8'b11001000;
	12'h0x501: q<=8'b10101001;
	12'h0x502: q<=8'b00000000;
	12'h0x503: q<=8'b10010001;
	12'h0x504: q<=8'b01110100;
	12'h0x505: q<=8'b11001000;
	12'h0x506: q<=8'b10010001;
	12'h0x507: q<=8'b01110100;
	12'h0x508: q<=8'b11001000;
	12'h0x509: q<=8'b10010001;
	12'h0x50a: q<=8'b01110100;
	12'h0x50b: q<=8'b10101001;
	12'h0x50c: q<=8'b10100000;
	12'h0x50d: q<=8'b11001000;
	12'h0x50e: q<=8'b10010001;
	12'h0x50f: q<=8'b01110100;
	12'h0x510: q<=8'b11001000;
	12'h0x511: q<=8'b10100101;
	12'h0x512: q<=8'b01100011;
	12'h0x513: q<=8'b01001001;
	12'h0x514: q<=8'b11111111;
	12'h0x515: q<=8'b00011000;
	12'h0x516: q<=8'b01101001;
	12'h0x517: q<=8'b00000001;
	12'h0x518: q<=8'b10010001;
	12'h0x519: q<=8'b01110100;
	12'h0x51a: q<=8'b11001000;
	12'h0x51b: q<=8'b10100101;
	12'h0x51c: q<=8'b01100100;
	12'h0x51d: q<=8'b01001001;
	12'h0x51e: q<=8'b11111111;
	12'h0x51f: q<=8'b01101001;
	12'h0x520: q<=8'b00000000;
	12'h0x521: q<=8'b00101001;
	12'h0x522: q<=8'b00011111;
	12'h0x523: q<=8'b10010001;
	12'h0x524: q<=8'b01110100;
	12'h0x525: q<=8'b11001000;
	12'h0x526: q<=8'b10100101;
	12'h0x527: q<=8'b01100001;
	12'h0x528: q<=8'b01001001;
	12'h0x529: q<=8'b11111111;
	12'h0x52a: q<=8'b00011000;
	12'h0x52b: q<=8'b01101001;
	12'h0x52c: q<=8'b00000001;
	12'h0x52d: q<=8'b10010001;
	12'h0x52e: q<=8'b01110100;
	12'h0x52f: q<=8'b11001000;
	12'h0x530: q<=8'b10100101;
	12'h0x531: q<=8'b01100010;
	12'h0x532: q<=8'b01001001;
	12'h0x533: q<=8'b11111111;
	12'h0x534: q<=8'b01101001;
	12'h0x535: q<=8'b00000000;
	12'h0x536: q<=8'b00101001;
	12'h0x537: q<=8'b00011111;
	12'h0x538: q<=8'b10010001;
	12'h0x539: q<=8'b01110100;
	12'h0x53a: q<=8'b11001000;
	12'h0x53b: q<=8'b11000000;
	12'h0x53c: q<=8'b11110000;
	12'h0x53d: q<=8'b10010000;
	12'h0x53e: q<=8'b00000110;
	12'h0x53f: q<=8'b10001000;
	12'h0x540: q<=8'b00100000;
	12'h0x541: q<=8'b01011111;
	12'h0x542: q<=8'b11011111;
	12'h0x543: q<=8'b10100000;
	12'h0x544: q<=8'b00000000;
	12'h0x545: q<=8'b11000110;
	12'h0x546: q<=8'b01010110;
	12'h0x547: q<=8'b00110000;
	12'h0x548: q<=8'b00000111;
	12'h0x549: q<=8'b11000110;
	12'h0x54a: q<=8'b00110111;
	12'h0x54b: q<=8'b00110000;
	12'h0x54c: q<=8'b00000011;
	12'h0x54d: q<=8'b01001100;
	12'h0x54e: q<=8'b10110000;
	12'h0x54f: q<=8'b10110100;
	12'h0x550: q<=8'b10011000;
	12'h0x551: q<=8'b11110000;
	12'h0x552: q<=8'b00000100;
	12'h0x553: q<=8'b10001000;
	12'h0x554: q<=8'b00100000;
	12'h0x555: q<=8'b01011111;
	12'h0x556: q<=8'b11011111;
	12'h0x557: q<=8'b10100101;
	12'h0x558: q<=8'b10110101;
	12'h0x559: q<=8'b11110000;
	12'h0x55a: q<=8'b00001010;
	12'h0x55b: q<=8'b10100101;
	12'h0x55c: q<=8'b01000110;
	12'h0x55d: q<=8'b11001001;
	12'h0x55e: q<=8'b00001010;
	12'h0x55f: q<=8'b10010000;
	12'h0x560: q<=8'b00000100;
	12'h0x561: q<=8'b10101001;
	12'h0x562: q<=8'b01111010;
	12'h0x563: q<=8'b10000101;
	12'h0x564: q<=8'b01010011;
	12'h0x565: q<=8'b10101001;
	12'h0x566: q<=8'b00000001;
	12'h0x567: q<=8'b01001100;
	12'h0x568: q<=8'b01101010;
	12'h0x569: q<=8'b11011111;
	12'h0x56a: q<=8'b01001000;
	12'h0x56b: q<=8'b10100000;
	12'h0x56c: q<=8'b00000000;
	12'h0x56d: q<=8'b10011000;
	12'h0x56e: q<=8'b10010001;
	12'h0x56f: q<=8'b01110100;
	12'h0x570: q<=8'b11001000;
	12'h0x571: q<=8'b10010001;
	12'h0x572: q<=8'b01110100;
	12'h0x573: q<=8'b11001000;
	12'h0x574: q<=8'b10010001;
	12'h0x575: q<=8'b01110100;
	12'h0x576: q<=8'b11001000;
	12'h0x577: q<=8'b01101000;
	12'h0x578: q<=8'b10010001;
	12'h0x579: q<=8'b01110100;
	12'h0x57a: q<=8'b10101001;
	12'h0x57b: q<=8'b00000100;
	12'h0x57c: q<=8'b00011000;
	12'h0x57d: q<=8'b01100101;
	12'h0x57e: q<=8'b01110100;
	12'h0x57f: q<=8'b10000101;
	12'h0x580: q<=8'b01110100;
	12'h0x581: q<=8'b10010000;
	12'h0x582: q<=8'b00000010;
	12'h0x583: q<=8'b11100110;
	12'h0x584: q<=8'b01110101;
	12'h0x585: q<=8'b01100000;
	12'h0x586: q<=8'b10101001;
	12'h0x587: q<=8'b00000001;
	12'h0x588: q<=8'b10000101;
	12'h0x589: q<=8'b10011110;
	12'h0x58a: q<=8'b10101101;
	12'h0x58b: q<=8'b00000010;
	12'h0x58c: q<=8'b00000010;
	12'h0x58d: q<=8'b11110000;
	12'h0x58e: q<=8'b00011101;
	12'h0x58f: q<=8'b11001001;
	12'h0x590: q<=8'b11110000;
	12'h0x591: q<=8'b10110000;
	12'h0x592: q<=8'b00011001;
	12'h0x593: q<=8'b10000101;
	12'h0x594: q<=8'b01010111;
	12'h0x595: q<=8'b10000101;
	12'h0x596: q<=8'b00101111;
	12'h0x597: q<=8'b10101101;
	12'h0x598: q<=8'b00000001;
	12'h0x599: q<=8'b00000010;
	12'h0x59a: q<=8'b11001001;
	12'h0x59b: q<=8'b10000001;
	12'h0x59c: q<=8'b11110000;
	12'h0x59d: q<=8'b00001110;
	12'h0x59e: q<=8'b10101100;
	12'h0x59f: q<=8'b00000000;
	12'h0x5a0: q<=8'b00000010;
	12'h0x5a1: q<=8'b10100101;
	12'h0x5a2: q<=8'b01010001;
	12'h0x5a3: q<=8'b01001010;
	12'h0x5a4: q<=8'b00101001;
	12'h0x5a5: q<=8'b00000111;
	12'h0x5a6: q<=8'b00011000;
	12'h0x5a7: q<=8'b01101001;
	12'h0x5a8: q<=8'b00000001;
	12'h0x5a9: q<=8'b00100000;
	12'h0x5aa: q<=8'b10100000;
	12'h0x5ab: q<=8'b10111101;
	12'h0x5ac: q<=8'b01100000;
	12'h0x5ad: q<=8'b10101101;
	12'h0x5ae: q<=8'b00000110;
	12'h0x5af: q<=8'b00000001;
	12'h0x5b0: q<=8'b00110000;
	12'h0x5b1: q<=8'b00100100;
	12'h0x5b2: q<=8'b10100010;
	12'h0x5b3: q<=8'b00000110;
	12'h0x5b4: q<=8'b10000110;
	12'h0x5b5: q<=8'b00110111;
	12'h0x5b6: q<=8'b10100110;
	12'h0x5b7: q<=8'b00110111;
	12'h0x5b8: q<=8'b10111101;
	12'h0x5b9: q<=8'b11011111;
	12'h0x5ba: q<=8'b00000010;
	12'h0x5bb: q<=8'b11110000;
	12'h0x5bc: q<=8'b00010101;
	12'h0x5bd: q<=8'b10000101;
	12'h0x5be: q<=8'b01010111;
	12'h0x5bf: q<=8'b10111101;
	12'h0x5c0: q<=8'b10000011;
	12'h0x5c1: q<=8'b00000010;
	12'h0x5c2: q<=8'b00101001;
	12'h0x5c3: q<=8'b00011000;
	12'h0x5c4: q<=8'b01001010;
	12'h0x5c5: q<=8'b01001010;
	12'h0x5c6: q<=8'b01001010;
	12'h0x5c7: q<=8'b10000101;
	12'h0x5c8: q<=8'b01010101;
	12'h0x5c9: q<=8'b10111101;
	12'h0x5ca: q<=8'b10000011;
	12'h0x5cb: q<=8'b00000010;
	12'h0x5cc: q<=8'b00101001;
	12'h0x5cd: q<=8'b00000111;
	12'h0x5ce: q<=8'b00001010;
	12'h0x5cf: q<=8'b00100000;
	12'h0x5d0: q<=8'b11010111;
	12'h0x5d1: q<=8'b10110101;
	12'h0x5d2: q<=8'b11000110;
	12'h0x5d3: q<=8'b00110111;
	12'h0x5d4: q<=8'b00010000;
	12'h0x5d5: q<=8'b11100000;
	12'h0x5d6: q<=8'b01100000;
	12'h0x5d7: q<=8'b10101000;
	12'h0x5d8: q<=8'b10111001;
	12'h0x5d9: q<=8'b11100010;
	12'h0x5da: q<=8'b10110101;
	12'h0x5db: q<=8'b01001000;
	12'h0x5dc: q<=8'b10111001;
	12'h0x5dd: q<=8'b11100001;
	12'h0x5de: q<=8'b10110101;
	12'h0x5df: q<=8'b01001000;
	12'h0x5e0: q<=8'b01100000;
	12'h0x5e1: q<=8'b11101010;
	12'h0x5e2: q<=8'b10110101;
	12'h0x5e3: q<=8'b00011010;
	12'h0x5e4: q<=8'b10110111;
	12'h0x5e5: q<=8'b00001110;
	12'h0x5e6: q<=8'b10110110;
	12'h0x5e7: q<=8'b00100001;
	12'h0x5e8: q<=8'b10110110;
	12'h0x5e9: q<=8'b10011010;
	12'h0x5ea: q<=8'b10110110;
	12'h0x5eb: q<=8'b10101001;
	12'h0x5ec: q<=8'b00000011;
	12'h0x5ed: q<=8'b10000101;
	12'h0x5ee: q<=8'b10011110;
	12'h0x5ef: q<=8'b10111101;
	12'h0x5f0: q<=8'b10000011;
	12'h0x5f1: q<=8'b00000010;
	12'h0x5f2: q<=8'b00110000;
	12'h0x5f3: q<=8'b00001110;
	12'h0x5f4: q<=8'b10111100;
	12'h0x5f5: q<=8'b10111001;
	12'h0x5f6: q<=8'b00000010;
	12'h0x5f7: q<=8'b10100110;
	12'h0x5f8: q<=8'b01010101;
	12'h0x5f9: q<=8'b10111101;
	12'h0x5fa: q<=8'b00001011;
	12'h0x5fb: q<=8'b10110110;
	12'h0x5fc: q<=8'b00100000;
	12'h0x5fd: q<=8'b10100000;
	12'h0x5fe: q<=8'b10111101;
	12'h0x5ff: q<=8'b10111000;
	12'h0x600: q<=8'b01010000;
	12'h0x601: q<=8'b00001000;
	12'h0x602: q<=8'b00100000;
	12'h0x603: q<=8'b00110100;
	12'h0x604: q<=8'b10110110;
	12'h0x605: q<=8'b10100000;
	12'h0x606: q<=8'b00000000;
	12'h0x607: q<=8'b00100000;
	12'h0x608: q<=8'b11001011;
	12'h0x609: q<=8'b10111101;
	12'h0x60a: q<=8'b01100000;
	12'h0x60b: q<=8'b00000000;
	12'h0x60c: q<=8'b00000000;
	12'h0x60d: q<=8'b00000000;
	12'h0x60e: q<=8'b00000000;
	12'h0x60f: q<=8'b10111101;
	12'h0x610: q<=8'b10001010;
	12'h0x611: q<=8'b00000010;
	12'h0x612: q<=8'b00101001;
	12'h0x613: q<=8'b00000011;
	12'h0x614: q<=8'b10101000;
	12'h0x615: q<=8'b10111001;
	12'h0x616: q<=8'b00011110;
	12'h0x617: q<=8'b10110110;
	12'h0x618: q<=8'b10111100;
	12'h0x619: q<=8'b10111001;
	12'h0x61a: q<=8'b00000010;
	12'h0x61b: q<=8'b01001100;
	12'h0x61c: q<=8'b11111101;
	12'h0x61d: q<=8'b10111100;
	12'h0x61e: q<=8'b00011010;
	12'h0x61f: q<=8'b00011010;
	12'h0x620: q<=8'b01001010;
	12'h0x621: q<=8'b01001100;
	12'h0x622: q<=8'b10111100;
	12'h0x623: q<=8'b10111001;
	12'h0x624: q<=8'b00000010;
	12'h0x625: q<=8'b10100101;
	12'h0x626: q<=8'b00000011;
	12'h0x627: q<=8'b00101001;
	12'h0x628: q<=8'b00000011;
	12'h0x629: q<=8'b00001010;
	12'h0x62a: q<=8'b00011000;
	12'h0x62b: q<=8'b01101001;
	12'h0x62c: q<=8'b00010010;
	12'h0x62d: q<=8'b01001100;
	12'h0x62e: q<=8'b11111101;
	12'h0x62f: q<=8'b10111100;
	12'h0x630: q<=8'b00010010;
	12'h0x631: q<=8'b00010100;
	12'h0x632: q<=8'b00010110;
	12'h0x633: q<=8'b00011000;
	12'h0x634: q<=8'b10100101;
	12'h0x635: q<=8'b01010111;
	12'h0x636: q<=8'b10000101;
	12'h0x637: q<=8'b00101111;
	12'h0x638: q<=8'b10111100;
	12'h0x639: q<=8'b10111001;
	12'h0x63a: q<=8'b00000010;
	12'h0x63b: q<=8'b10111001;
	12'h0x63c: q<=8'b11001110;
	12'h0x63d: q<=8'b00000011;
	12'h0x63e: q<=8'b10000101;
	12'h0x63f: q<=8'b01010110;
	12'h0x640: q<=8'b10111001;
	12'h0x641: q<=8'b11011110;
	12'h0x642: q<=8'b00000011;
	12'h0x643: q<=8'b10000101;
	12'h0x644: q<=8'b01011000;
	12'h0x645: q<=8'b10111101;
	12'h0x646: q<=8'b11001100;
	12'h0x647: q<=8'b00000010;
	12'h0x648: q<=8'b00101001;
	12'h0x649: q<=8'b00001111;
	12'h0x64a: q<=8'b10101000;
	12'h0x64b: q<=8'b10100101;
	12'h0x64c: q<=8'b01010110;
	12'h0x64d: q<=8'b01001001;
	12'h0x64e: q<=8'b10000000;
	12'h0x64f: q<=8'b00011000;
	12'h0x650: q<=8'b01111001;
	12'h0x651: q<=8'b10001011;
	12'h0x652: q<=8'b10110110;
	12'h0x653: q<=8'b01010000;
	12'h0x654: q<=8'b00001001;
	12'h0x655: q<=8'b00010000;
	12'h0x656: q<=8'b00000101;
	12'h0x657: q<=8'b10101001;
	12'h0x658: q<=8'b01111111;
	12'h0x659: q<=8'b10111000;
	12'h0x65a: q<=8'b01010000;
	12'h0x65b: q<=8'b00000010;
	12'h0x65c: q<=8'b10101001;
	12'h0x65d: q<=8'b10000000;
	12'h0x65e: q<=8'b01001001;
	12'h0x65f: q<=8'b10000000;
	12'h0x660: q<=8'b10000101;
	12'h0x661: q<=8'b00101110;
	12'h0x662: q<=8'b10100101;
	12'h0x663: q<=8'b01011000;
	12'h0x664: q<=8'b01001001;
	12'h0x665: q<=8'b10000000;
	12'h0x666: q<=8'b00011000;
	12'h0x667: q<=8'b01111001;
	12'h0x668: q<=8'b10000111;
	12'h0x669: q<=8'b10110110;
	12'h0x66a: q<=8'b01010000;
	12'h0x66b: q<=8'b00001001;
	12'h0x66c: q<=8'b00010000;
	12'h0x66d: q<=8'b00000101;
	12'h0x66e: q<=8'b10101001;
	12'h0x66f: q<=8'b01111111;
	12'h0x670: q<=8'b10111000;
	12'h0x671: q<=8'b01010000;
	12'h0x672: q<=8'b00000010;
	12'h0x673: q<=8'b10101001;
	12'h0x674: q<=8'b10000000;
	12'h0x675: q<=8'b01001001;
	12'h0x676: q<=8'b10000000;
	12'h0x677: q<=8'b10000101;
	12'h0x678: q<=8'b00110000;
	12'h0x679: q<=8'b10101100;
	12'h0x67a: q<=8'b00010010;
	12'h0x67b: q<=8'b00000001;
	12'h0x67c: q<=8'b10111001;
	12'h0x67d: q<=8'b11011100;
	12'h0x67e: q<=8'b10111100;
	12'h0x67f: q<=8'b10000101;
	12'h0x680: q<=8'b01011001;
	12'h0x681: q<=8'b10111001;
	12'h0x682: q<=8'b11101100;
	12'h0x683: q<=8'b10111100;
	12'h0x684: q<=8'b10000101;
	12'h0x685: q<=8'b01011010;
	12'h0x686: q<=8'b01100000;
	12'h0x687: q<=8'b00000000;
	12'h0x688: q<=8'b00010000;
	12'h0x689: q<=8'b00011111;
	12'h0x68a: q<=8'b00101000;
	12'h0x68b: q<=8'b00101100;
	12'h0x68c: q<=8'b00101000;
	12'h0x68d: q<=8'b00011111;
	12'h0x68e: q<=8'b00010000;
	12'h0x68f: q<=8'b00000000;
	12'h0x690: q<=8'b11110000;
	12'h0x691: q<=8'b11100001;
	12'h0x692: q<=8'b11011000;
	12'h0x693: q<=8'b11010100;
	12'h0x694: q<=8'b11011000;
	12'h0x695: q<=8'b11100001;
	12'h0x696: q<=8'b11110000;
	12'h0x697: q<=8'b00000000;
	12'h0x698: q<=8'b00010000;
	12'h0x699: q<=8'b00011111;
	12'h0x69a: q<=8'b00101000;
	12'h0x69b: q<=8'b10111101;
	12'h0x69c: q<=8'b11011111;
	12'h0x69d: q<=8'b00000010;
	12'h0x69e: q<=8'b10000101;
	12'h0x69f: q<=8'b01010111;
	12'h0x6a0: q<=8'b10111100;
	12'h0x6a1: q<=8'b10111001;
	12'h0x6a2: q<=8'b00000010;
	12'h0x6a3: q<=8'b10111001;
	12'h0x6a4: q<=8'b11001110;
	12'h0x6a5: q<=8'b00000011;
	12'h0x6a6: q<=8'b10000101;
	12'h0x6a7: q<=8'b01010110;
	12'h0x6a8: q<=8'b10111001;
	12'h0x6a9: q<=8'b11011110;
	12'h0x6aa: q<=8'b00000011;
	12'h0x6ab: q<=8'b10000101;
	12'h0x6ac: q<=8'b01011000;
	12'h0x6ad: q<=8'b10111101;
	12'h0x6ae: q<=8'b11001100;
	12'h0x6af: q<=8'b00000010;
	12'h0x6b0: q<=8'b00010000;
	12'h0x6b1: q<=8'b00100011;
	12'h0x6b2: q<=8'b10011000;
	12'h0x6b3: q<=8'b00011000;
	12'h0x6b4: q<=8'b01101001;
	12'h0x6b5: q<=8'b00000001;
	12'h0x6b6: q<=8'b00101001;
	12'h0x6b7: q<=8'b00001111;
	12'h0x6b8: q<=8'b10101000;
	12'h0x6b9: q<=8'b10111001;
	12'h0x6ba: q<=8'b11001110;
	12'h0x6bb: q<=8'b00000011;
	12'h0x6bc: q<=8'b00111000;
	12'h0x6bd: q<=8'b11100101;
	12'h0x6be: q<=8'b01010110;
	12'h0x6bf: q<=8'b00100000;
	12'h0x6c0: q<=8'b11111010;
	12'h0x6c1: q<=8'b10110110;
	12'h0x6c2: q<=8'b00011000;
	12'h0x6c3: q<=8'b01100101;
	12'h0x6c4: q<=8'b01010110;
	12'h0x6c5: q<=8'b10000101;
	12'h0x6c6: q<=8'b01010110;
	12'h0x6c7: q<=8'b10111001;
	12'h0x6c8: q<=8'b11011110;
	12'h0x6c9: q<=8'b00000011;
	12'h0x6ca: q<=8'b00111000;
	12'h0x6cb: q<=8'b11100101;
	12'h0x6cc: q<=8'b01011000;
	12'h0x6cd: q<=8'b00100000;
	12'h0x6ce: q<=8'b11111010;
	12'h0x6cf: q<=8'b10110110;
	12'h0x6d0: q<=8'b00011000;
	12'h0x6d1: q<=8'b01100101;
	12'h0x6d2: q<=8'b01011000;
	12'h0x6d3: q<=8'b10000101;
	12'h0x6d4: q<=8'b01011000;
	12'h0x6d5: q<=8'b00100000;
	12'h0x6d6: q<=8'b10011000;
	12'h0x6d7: q<=8'b11000000;
	12'h0x6d8: q<=8'b10100010;
	12'h0x6d9: q<=8'b01100001;
	12'h0x6da: q<=8'b00100000;
	12'h0x6db: q<=8'b01100101;
	12'h0x6dc: q<=8'b11000111;
	12'h0x6dd: q<=8'b10101001;
	12'h0x6de: q<=8'b00000000;
	12'h0x6df: q<=8'b10000101;
	12'h0x6e0: q<=8'b10101001;
	12'h0x6e1: q<=8'b00100000;
	12'h0x6e2: q<=8'b00111110;
	12'h0x6e3: q<=8'b10111101;
	12'h0x6e4: q<=8'b10000100;
	12'h0x6e5: q<=8'b10101001;
	12'h0x6e6: q<=8'b10100101;
	12'h0x6e7: q<=8'b00000011;
	12'h0x6e8: q<=8'b00101001;
	12'h0x6e9: q<=8'b00000011;
	12'h0x6ea: q<=8'b00001010;
	12'h0x6eb: q<=8'b00011000;
	12'h0x6ec: q<=8'b01101001;
	12'h0x6ed: q<=8'b01001110;
	12'h0x6ee: q<=8'b10101000;
	12'h0x6ef: q<=8'b10111110;
	12'h0x6f0: q<=8'b11001001;
	12'h0x6f1: q<=8'b11001110;
	12'h0x6f2: q<=8'b10111001;
	12'h0x6f3: q<=8'b11001000;
	12'h0x6f4: q<=8'b11001110;
	12'h0x6f5: q<=8'b10100100;
	12'h0x6f6: q<=8'b10101001;
	12'h0x6f7: q<=8'b01001100;
	12'h0x6f8: q<=8'b01011001;
	12'h0x6f9: q<=8'b11011111;
	12'h0x6fa: q<=8'b10000101;
	12'h0x6fb: q<=8'b00101001;
	12'h0x6fc: q<=8'b10111101;
	12'h0x6fd: q<=8'b11001100;
	12'h0x6fe: q<=8'b00000010;
	12'h0x6ff: q<=8'b00101001;
	12'h0x700: q<=8'b00000111;
	12'h0x701: q<=8'b10000101;
	12'h0x702: q<=8'b00101100;
	12'h0x703: q<=8'b10000110;
	12'h0x704: q<=8'b00101011;
	12'h0x705: q<=8'b10100010;
	12'h0x706: q<=8'b00000010;
	12'h0x707: q<=8'b10101001;
	12'h0x708: q<=8'b00000000;
	12'h0x709: q<=8'b01000110;
	12'h0x70a: q<=8'b00101100;
	12'h0x70b: q<=8'b10010000;
	12'h0x70c: q<=8'b00000011;
	12'h0x70d: q<=8'b00011000;
	12'h0x70e: q<=8'b01100101;
	12'h0x70f: q<=8'b00101001;
	12'h0x710: q<=8'b00001010;
	12'h0x711: q<=8'b00001000;
	12'h0x712: q<=8'b01101010;
	12'h0x713: q<=8'b00101000;
	12'h0x714: q<=8'b01101010;
	12'h0x715: q<=8'b11001010;
	12'h0x716: q<=8'b00010000;
	12'h0x717: q<=8'b11110001;
	12'h0x718: q<=8'b10100110;
	12'h0x719: q<=8'b00101011;
	12'h0x71a: q<=8'b01100000;
	12'h0x71b: q<=8'b10101001;
	12'h0x71c: q<=8'b00000100;
	12'h0x71d: q<=8'b10101100;
	12'h0x71e: q<=8'b01001000;
	12'h0x71f: q<=8'b00000001;
	12'h0x720: q<=8'b00110000;
	12'h0x721: q<=8'b00000010;
	12'h0x722: q<=8'b10101001;
	12'h0x723: q<=8'b00000000;
	12'h0x724: q<=8'b10000101;
	12'h0x725: q<=8'b10011110;
	12'h0x726: q<=8'b10101101;
	12'h0x727: q<=8'b01001000;
	12'h0x728: q<=8'b00000001;
	12'h0x729: q<=8'b00011000;
	12'h0x72a: q<=8'b01101001;
	12'h0x72b: q<=8'b01000000;
	12'h0x72c: q<=8'b01001010;
	12'h0x72d: q<=8'b01001010;
	12'h0x72e: q<=8'b01001010;
	12'h0x72f: q<=8'b01001010;
	12'h0x730: q<=8'b11001001;
	12'h0x731: q<=8'b00000101;
	12'h0x732: q<=8'b10010000;
	12'h0x733: q<=8'b00000010;
	12'h0x734: q<=8'b10101001;
	12'h0x735: q<=8'b00000000;
	12'h0x736: q<=8'b10101000;
	12'h0x737: q<=8'b10111001;
	12'h0x738: q<=8'b01010101;
	12'h0x739: q<=8'b10110111;
	12'h0x73a: q<=8'b10000101;
	12'h0x73b: q<=8'b00101001;
	12'h0x73c: q<=8'b10111101;
	12'h0x73d: q<=8'b10000011;
	12'h0x73e: q<=8'b00000010;
	12'h0x73f: q<=8'b00110000;
	12'h0x740: q<=8'b00001011;
	12'h0x741: q<=8'b10111100;
	12'h0x742: q<=8'b10111001;
	12'h0x743: q<=8'b00000010;
	12'h0x744: q<=8'b10100101;
	12'h0x745: q<=8'b00101001;
	12'h0x746: q<=8'b00100000;
	12'h0x747: q<=8'b10100000;
	12'h0x748: q<=8'b10111101;
	12'h0x749: q<=8'b10111000;
	12'h0x74a: q<=8'b01010000;
	12'h0x74b: q<=8'b00001000;
	12'h0x74c: q<=8'b00100000;
	12'h0x74d: q<=8'b00110100;
	12'h0x74e: q<=8'b10110110;
	12'h0x74f: q<=8'b10100100;
	12'h0x750: q<=8'b00101001;
	12'h0x751: q<=8'b00100000;
	12'h0x752: q<=8'b11001011;
	12'h0x753: q<=8'b10111101;
	12'h0x754: q<=8'b01100000;
	12'h0x755: q<=8'b00001101;
	12'h0x756: q<=8'b00001100;
	12'h0x757: q<=8'b00001011;
	12'h0x758: q<=8'b00001010;
	12'h0x759: q<=8'b00001001;
	12'h0x75a: q<=8'b00001001;
	12'h0x75b: q<=8'b10100010;
	12'h0x75c: q<=8'b00001011;
	12'h0x75d: q<=8'b10000110;
	12'h0x75e: q<=8'b00110111;
	12'h0x75f: q<=8'b10100110;
	12'h0x760: q<=8'b00110111;
	12'h0x761: q<=8'b10111101;
	12'h0x762: q<=8'b11010011;
	12'h0x763: q<=8'b00000010;
	12'h0x764: q<=8'b11110000;
	12'h0x765: q<=8'b00011011;
	12'h0x766: q<=8'b10000101;
	12'h0x767: q<=8'b01010111;
	12'h0x768: q<=8'b10000101;
	12'h0x769: q<=8'b00101111;
	12'h0x76a: q<=8'b11100000;
	12'h0x76b: q<=8'b00001000;
	12'h0x76c: q<=8'b10111100;
	12'h0x76d: q<=8'b10101101;
	12'h0x76e: q<=8'b00000010;
	12'h0x76f: q<=8'b10110000;
	12'h0x770: q<=8'b00000101;
	12'h0x771: q<=8'b10101001;
	12'h0x772: q<=8'b00001000;
	12'h0x773: q<=8'b10111000;
	12'h0x774: q<=8'b01010000;
	12'h0x775: q<=8'b00001000;
	12'h0x776: q<=8'b10100101;
	12'h0x777: q<=8'b00000011;
	12'h0x778: q<=8'b00001010;
	12'h0x779: q<=8'b00101001;
	12'h0x77a: q<=8'b00000110;
	12'h0x77b: q<=8'b00011000;
	12'h0x77c: q<=8'b01101001;
	12'h0x77d: q<=8'b00100000;
	12'h0x77e: q<=8'b00100000;
	12'h0x77f: q<=8'b11111101;
	12'h0x780: q<=8'b10111100;
	12'h0x781: q<=8'b11000110;
	12'h0x782: q<=8'b00110111;
	12'h0x783: q<=8'b00010000;
	12'h0x784: q<=8'b11011010;
	12'h0x785: q<=8'b10100000;
	12'h0x786: q<=8'b00000100;
	12'h0x787: q<=8'b10101101;
	12'h0x788: q<=8'b00110101;
	12'h0x789: q<=8'b00000001;
	12'h0x78a: q<=8'b11001001;
	12'h0x78b: q<=8'b00000110;
	12'h0x78c: q<=8'b10010000;
	12'h0x78d: q<=8'b00001000;
	12'h0x78e: q<=8'b10100000;
	12'h0x78f: q<=8'b00001011;
	12'h0x790: q<=8'b11001001;
	12'h0x791: q<=8'b00001000;
	12'h0x792: q<=8'b10010000;
	12'h0x793: q<=8'b00000010;
	12'h0x794: q<=8'b10100000;
	12'h0x795: q<=8'b00001100;
	12'h0x796: q<=8'b10001100;
	12'h0x797: q<=8'b00001000;
	12'h0x798: q<=8'b00001000;
	12'h0x799: q<=8'b01100000;
	12'h0x79a: q<=8'b10100000;
	12'h0x79b: q<=8'b00000000;
	12'h0x79c: q<=8'b10000100;
	12'h0x79d: q<=8'b10011110;
	12'h0x79e: q<=8'b10100010;
	12'h0x79f: q<=8'b00000111;
	12'h0x7a0: q<=8'b10000110;
	12'h0x7a1: q<=8'b00110111;
	12'h0x7a2: q<=8'b10100110;
	12'h0x7a3: q<=8'b00110111;
	12'h0x7a4: q<=8'b10111101;
	12'h0x7a5: q<=8'b00001010;
	12'h0x7a6: q<=8'b00000011;
	12'h0x7a7: q<=8'b11110000;
	12'h0x7a8: q<=8'b00101001;
	12'h0x7a9: q<=8'b10000101;
	12'h0x7aa: q<=8'b01010111;
	12'h0x7ab: q<=8'b10111101;
	12'h0x7ac: q<=8'b11111010;
	12'h0x7ad: q<=8'b00000010;
	12'h0x7ae: q<=8'b10000101;
	12'h0x7af: q<=8'b00101001;
	12'h0x7b0: q<=8'b10111100;
	12'h0x7b1: q<=8'b00000010;
	12'h0x7b2: q<=8'b00000011;
	12'h0x7b3: q<=8'b11000000;
	12'h0x7b4: q<=8'b00000001;
	12'h0x7b5: q<=8'b11010000;
	12'h0x7b6: q<=8'b00000110;
	12'h0x7b7: q<=8'b00100000;
	12'h0x7b8: q<=8'b11101011;
	12'h0x7b9: q<=8'b10110111;
	12'h0x7ba: q<=8'b10111000;
	12'h0x7bb: q<=8'b01010000;
	12'h0x7bc: q<=8'b00010101;
	12'h0x7bd: q<=8'b10111101;
	12'h0x7be: q<=8'b00010010;
	12'h0x7bf: q<=8'b00000011;
	12'h0x7c0: q<=8'b01001010;
	12'h0x7c1: q<=8'b00101001;
	12'h0x7c2: q<=8'b11111110;
	12'h0x7c3: q<=8'b11000000;
	12'h0x7c4: q<=8'b00000010;
	12'h0x7c5: q<=8'b10010000;
	12'h0x7c6: q<=8'b00000010;
	12'h0x7c7: q<=8'b10101001;
	12'h0x7c8: q<=8'b00000000;
	12'h0x7c9: q<=8'b00011000;
	12'h0x7ca: q<=8'b01111001;
	12'h0x7cb: q<=8'b11100101;
	12'h0x7cc: q<=8'b10110111;
	12'h0x7cd: q<=8'b10100100;
	12'h0x7ce: q<=8'b00101001;
	12'h0x7cf: q<=8'b00100000;
	12'h0x7d0: q<=8'b11111101;
	12'h0x7d1: q<=8'b10111100;
	12'h0x7d2: q<=8'b11000110;
	12'h0x7d3: q<=8'b00110111;
	12'h0x7d4: q<=8'b00010000;
	12'h0x7d5: q<=8'b11001100;
	12'h0x7d6: q<=8'b10101101;
	12'h0x7d7: q<=8'b00100000;
	12'h0x7d8: q<=8'b00000111;
	12'h0x7d9: q<=8'b11110000;
	12'h0x7da: q<=8'b00001001;
	12'h0x7db: q<=8'b10100101;
	12'h0x7dc: q<=8'b10011111;
	12'h0x7dd: q<=8'b11001001;
	12'h0x7de: q<=8'b00001101;
	12'h0x7df: q<=8'b10010000;
	12'h0x7e0: q<=8'b00000011;
	12'h0x7e1: q<=8'b10001101;
	12'h0x7e2: q<=8'b11111111;
	12'h0x7e3: q<=8'b00000001;
	12'h0x7e4: q<=8'b01100000;
	12'h0x7e5: q<=8'b00000000;
	12'h0x7e6: q<=8'b00000000;
	12'h0x7e7: q<=8'b01011010;
	12'h0x7e8: q<=8'b01011000;
	12'h0x7e9: q<=8'b01010110;
	12'h0x7ea: q<=8'b00011100;
	12'h0x7eb: q<=8'b10100100;
	12'h0x7ec: q<=8'b00101001;
	12'h0x7ed: q<=8'b10111001;
	12'h0x7ee: q<=8'b00110101;
	12'h0x7ef: q<=8'b00000100;
	12'h0x7f0: q<=8'b10000101;
	12'h0x7f1: q<=8'b01010110;
	12'h0x7f2: q<=8'b10111001;
	12'h0x7f3: q<=8'b01000101;
	12'h0x7f4: q<=8'b00000100;
	12'h0x7f5: q<=8'b10000101;
	12'h0x7f6: q<=8'b01011000;
	12'h0x7f7: q<=8'b00100000;
	12'h0x7f8: q<=8'b10011000;
	12'h0x7f9: q<=8'b11000000;
	12'h0x7fa: q<=8'b10100010;
	12'h0x7fb: q<=8'b01100001;
	12'h0x7fc: q<=8'b00100000;
	12'h0x7fd: q<=8'b01100101;
	12'h0x7fe: q<=8'b11000111;
	12'h0x7ff: q<=8'b10101110;
	12'h0x800: q<=8'b00111011;
	12'h0x801: q<=8'b00000001;
	12'h0x802: q<=8'b11001110;
	12'h0x803: q<=8'b00111100;
	12'h0x804: q<=8'b00000001;
	12'h0x805: q<=8'b11010000;
	12'h0x806: q<=8'b00001010;
	12'h0x807: q<=8'b11101000;
	12'h0x808: q<=8'b10001110;
	12'h0x809: q<=8'b00111011;
	12'h0x80a: q<=8'b00000001;
	12'h0x80b: q<=8'b10111101;
	12'h0x80c: q<=8'b00101010;
	12'h0x80d: q<=8'b10111000;
	12'h0x80e: q<=8'b10001101;
	12'h0x80f: q<=8'b00111100;
	12'h0x810: q<=8'b00000001;
	12'h0x811: q<=8'b10111100;
	12'h0x812: q<=8'b00111101;
	12'h0x813: q<=8'b10111000;
	12'h0x814: q<=8'b00110000;
	12'h0x815: q<=8'b00000011;
	12'h0x816: q<=8'b00100000;
	12'h0x817: q<=8'b01001110;
	12'h0x818: q<=8'b10111000;
	12'h0x819: q<=8'b10101101;
	12'h0x81a: q<=8'b00111011;
	12'h0x81b: q<=8'b00000001;
	12'h0x81c: q<=8'b00001010;
	12'h0x81d: q<=8'b00011000;
	12'h0x81e: q<=8'b01101001;
	12'h0x81f: q<=8'b00101000;
	12'h0x820: q<=8'b10101000;
	12'h0x821: q<=8'b10111110;
	12'h0x822: q<=8'b11001001;
	12'h0x823: q<=8'b11001110;
	12'h0x824: q<=8'b10111001;
	12'h0x825: q<=8'b11001000;
	12'h0x826: q<=8'b11001110;
	12'h0x827: q<=8'b01001100;
	12'h0x828: q<=8'b01010111;
	12'h0x829: q<=8'b11011111;
	12'h0x82a: q<=8'b00000010;
	12'h0x82b: q<=8'b00000010;
	12'h0x82c: q<=8'b00000010;
	12'h0x82d: q<=8'b00000010;
	12'h0x82e: q<=8'b00000010;
	12'h0x82f: q<=8'b00000100;
	12'h0x830: q<=8'b00000011;
	12'h0x831: q<=8'b00000010;
	12'h0x832: q<=8'b00000001;
	12'h0x833: q<=8'b00100000;
	12'h0x834: q<=8'b00000011;
	12'h0x835: q<=8'b00000011;
	12'h0x836: q<=8'b00000011;
	12'h0x837: q<=8'b00000011;
	12'h0x838: q<=8'b00000011;
	12'h0x839: q<=8'b00000011;
	12'h0x83a: q<=8'b00000011;
	12'h0x83b: q<=8'b00111011;
	12'h0x83c: q<=8'b10111000;
	12'h0x83d: q<=8'b00000000;
	12'h0x83e: q<=8'b00000010;
	12'h0x83f: q<=8'b00000010;
	12'h0x840: q<=8'b00000010;
	12'h0x841: q<=8'b00000010;
	12'h0x842: q<=8'b00000010;
	12'h0x843: q<=8'b00000010;
	12'h0x844: q<=8'b00000010;
	12'h0x845: q<=8'b00000100;
	12'h0x846: q<=8'b00000110;
	12'h0x847: q<=8'b11111111;
	12'h0x848: q<=8'b11111111;
	12'h0x849: q<=8'b11111111;
	12'h0x84a: q<=8'b11111111;
	12'h0x84b: q<=8'b11111111;
	12'h0x84c: q<=8'b11111111;
	12'h0x84d: q<=8'b11111111;
	12'h0x84e: q<=8'b10111001;
	12'h0x84f: q<=8'b01011000;
	12'h0x850: q<=8'b10111000;
	12'h0x851: q<=8'b01001000;
	12'h0x852: q<=8'b10111001;
	12'h0x853: q<=8'b01010111;
	12'h0x854: q<=8'b10111000;
	12'h0x855: q<=8'b01001000;
	12'h0x856: q<=8'b01100000;
	12'h0x857: q<=8'b01011110;
	12'h0x858: q<=8'b10111000;
	12'h0x859: q<=8'b01110100;
	12'h0x85a: q<=8'b10111000;
	12'h0x85b: q<=8'b10000111;
	12'h0x85c: q<=8'b10111000;
	12'h0x85d: q<=8'b10010101;
	12'h0x85e: q<=8'b10111000;
	12'h0x85f: q<=8'b10101001;
	12'h0x860: q<=8'b00001100;
	12'h0x861: q<=8'b10001101;
	12'h0x862: q<=8'b00001011;
	12'h0x863: q<=8'b00001000;
	12'h0x864: q<=8'b10000101;
	12'h0x865: q<=8'b00100100;
	12'h0x866: q<=8'b10101001;
	12'h0x867: q<=8'b00000100;
	12'h0x868: q<=8'b10001101;
	12'h0x869: q<=8'b00001010;
	12'h0x86a: q<=8'b00001000;
	12'h0x86b: q<=8'b10000101;
	12'h0x86c: q<=8'b00100011;
	12'h0x86d: q<=8'b10101001;
	12'h0x86e: q<=8'b00000000;
	12'h0x86f: q<=8'b10000101;
	12'h0x870: q<=8'b00100010;
	12'h0x871: q<=8'b10001101;
	12'h0x872: q<=8'b00001001;
	12'h0x873: q<=8'b00001000;
	12'h0x874: q<=8'b01100000;
	12'h0x875: q<=8'b10100100;
	12'h0x876: q<=8'b00100010;
	12'h0x877: q<=8'b10100010;
	12'h0x878: q<=8'b00000010;
	12'h0x879: q<=8'b10110101;
	12'h0x87a: q<=8'b00100010;
	12'h0x87b: q<=8'b01001000;
	12'h0x87c: q<=8'b10010100;
	12'h0x87d: q<=8'b00100010;
	12'h0x87e: q<=8'b10011000;
	12'h0x87f: q<=8'b10011101;
	12'h0x880: q<=8'b00001001;
	12'h0x881: q<=8'b00001000;
	12'h0x882: q<=8'b01101000;
	12'h0x883: q<=8'b10101000;
	12'h0x884: q<=8'b11001010;
	12'h0x885: q<=8'b00010000;
	12'h0x886: q<=8'b11110010;
	12'h0x887: q<=8'b01100000;
	12'h0x888: q<=8'b00100000;
	12'h0x889: q<=8'b10010110;
	12'h0x88a: q<=8'b11000001;
	12'h0x88b: q<=8'b10101001;
	12'h0x88c: q<=8'b01111111;
	12'h0x88d: q<=8'b10001101;
	12'h0x88e: q<=8'b00111001;
	12'h0x88f: q<=8'b00000001;
	12'h0x890: q<=8'b10101001;
	12'h0x891: q<=8'b00000100;
	12'h0x892: q<=8'b10001101;
	12'h0x893: q<=8'b00111010;
	12'h0x894: q<=8'b00000001;
	12'h0x895: q<=8'b01100000;
	12'h0x896: q<=8'b10101101;
	12'h0x897: q<=8'b00111001;
	12'h0x898: q<=8'b00000001;
	12'h0x899: q<=8'b10001101;
	12'h0x89a: q<=8'b11111100;
	12'h0x89b: q<=8'b00101111;
	12'h0x89c: q<=8'b10101101;
	12'h0x89d: q<=8'b00111010;
	12'h0x89e: q<=8'b00000001;
	12'h0x89f: q<=8'b00001001;
	12'h0x8a0: q<=8'b01110000;
	12'h0x8a1: q<=8'b10001101;
	12'h0x8a2: q<=8'b11111101;
	12'h0x8a3: q<=8'b00101111;
	12'h0x8a4: q<=8'b10101001;
	12'h0x8a5: q<=8'b11000000;
	12'h0x8a6: q<=8'b10001101;
	12'h0x8a7: q<=8'b11111111;
	12'h0x8a8: q<=8'b00101111;
	12'h0x8a9: q<=8'b10101101;
	12'h0x8aa: q<=8'b00111001;
	12'h0x8ab: q<=8'b00000001;
	12'h0x8ac: q<=8'b00111000;
	12'h0x8ad: q<=8'b11101001;
	12'h0x8ae: q<=8'b00100000;
	12'h0x8af: q<=8'b00010000;
	12'h0x8b0: q<=8'b00000101;
	12'h0x8b1: q<=8'b00101001;
	12'h0x8b2: q<=8'b01111111;
	12'h0x8b3: q<=8'b11001110;
	12'h0x8b4: q<=8'b00111010;
	12'h0x8b5: q<=8'b00000001;
	12'h0x8b6: q<=8'b10001101;
	12'h0x8b7: q<=8'b00111001;
	12'h0x8b8: q<=8'b00000001;
	12'h0x8b9: q<=8'b01100000;
	12'h0x8ba: q<=8'b10101001;
	12'h0x8bb: q<=8'b00111111;
	12'h0x8bc: q<=8'b10100010;
	12'h0x8bd: q<=8'b11110010;
	12'h0x8be: q<=8'b00100000;
	12'h0x8bf: q<=8'b00111001;
	12'h0x8c0: q<=8'b11011111;
	12'h0x8c1: q<=8'b10101001;
	12'h0x8c2: q<=8'b00000000;
	12'h0x8c3: q<=8'b10000101;
	12'h0x8c4: q<=8'b01101010;
	12'h0x8c5: q<=8'b10000101;
	12'h0x8c6: q<=8'b01101011;
	12'h0x8c7: q<=8'b10000101;
	12'h0x8c8: q<=8'b01101100;
	12'h0x8c9: q<=8'b10000101;
	12'h0x8ca: q<=8'b01101101;
	12'h0x8cb: q<=8'b10001101;
	12'h0x8cc: q<=8'b00000010;
	12'h0x8cd: q<=8'b00000010;
	12'h0x8ce: q<=8'b10000101;
	12'h0x8cf: q<=8'b01101000;
	12'h0x8d0: q<=8'b10000101;
	12'h0x8d1: q<=8'b01101001;
	12'h0x8d2: q<=8'b10101001;
	12'h0x8d3: q<=8'b11100000;
	12'h0x8d4: q<=8'b10000101;
	12'h0x8d5: q<=8'b01011111;
	12'h0x8d6: q<=8'b10101001;
	12'h0x8d7: q<=8'b11111111;
	12'h0x8d8: q<=8'b10000101;
	12'h0x8d9: q<=8'b01011011;
	12'h0x8da: q<=8'b00100000;
	12'h0x8db: q<=8'b01100111;
	12'h0x8dc: q<=8'b10111001;
	12'h0x8dd: q<=8'b10000101;
	12'h0x8de: q<=8'b01110111;
	12'h0x8df: q<=8'b10000110;
	12'h0x8e0: q<=8'b01110110;
	12'h0x8e1: q<=8'b10100010;
	12'h0x8e2: q<=8'b00001111;
	12'h0x8e3: q<=8'b10000110;
	12'h0x8e4: q<=8'b00110111;
	12'h0x8e5: q<=8'b10100110;
	12'h0x8e6: q<=8'b00110111;
	12'h0x8e7: q<=8'b10111101;
	12'h0x8e8: q<=8'b10000011;
	12'h0x8e9: q<=8'b00000010;
	12'h0x8ea: q<=8'b11110000;
	12'h0x8eb: q<=8'b01001001;
	12'h0x8ec: q<=8'b10000101;
	12'h0x8ed: q<=8'b01010111;
	12'h0x8ee: q<=8'b10111101;
	12'h0x8ef: q<=8'b01100011;
	12'h0x8f0: q<=8'b00000010;
	12'h0x8f1: q<=8'b10000101;
	12'h0x8f2: q<=8'b01010110;
	12'h0x8f3: q<=8'b10111101;
	12'h0x8f4: q<=8'b10100011;
	12'h0x8f5: q<=8'b00000010;
	12'h0x8f6: q<=8'b10000101;
	12'h0x8f7: q<=8'b01011000;
	12'h0x8f8: q<=8'b00100000;
	12'h0x8f9: q<=8'b10011000;
	12'h0x8fa: q<=8'b11000000;
	12'h0x8fb: q<=8'b10101001;
	12'h0x8fc: q<=8'b00000000;
	12'h0x8fd: q<=8'b10000101;
	12'h0x8fe: q<=8'b01110011;
	12'h0x8ff: q<=8'b00100000;
	12'h0x900: q<=8'b01000100;
	12'h0x901: q<=8'b10111001;
	12'h0x902: q<=8'b00100000;
	12'h0x903: q<=8'b10111010;
	12'h0x904: q<=8'b11000011;
	12'h0x905: q<=8'b10101001;
	12'h0x906: q<=8'b10100000;
	12'h0x907: q<=8'b00100000;
	12'h0x908: q<=8'b01101010;
	12'h0x909: q<=8'b10110101;
	12'h0x90a: q<=8'b00100000;
	12'h0x90b: q<=8'b01000100;
	12'h0x90c: q<=8'b10111001;
	12'h0x90d: q<=8'b10100010;
	12'h0x90e: q<=8'b01100001;
	12'h0x90f: q<=8'b00100000;
	12'h0x910: q<=8'b01110010;
	12'h0x911: q<=8'b11000111;
	12'h0x912: q<=8'b00100000;
	12'h0x913: q<=8'b01010101;
	12'h0x914: q<=8'b10111001;
	12'h0x915: q<=8'b00100000;
	12'h0x916: q<=8'b01101100;
	12'h0x917: q<=8'b11011111;
	12'h0x918: q<=8'b10100101;
	12'h0x919: q<=8'b00110111;
	12'h0x91a: q<=8'b00101001;
	12'h0x91b: q<=8'b00000111;
	12'h0x91c: q<=8'b11001001;
	12'h0x91d: q<=8'b00000111;
	12'h0x91e: q<=8'b11010000;
	12'h0x91f: q<=8'b00000010;
	12'h0x920: q<=8'b10101001;
	12'h0x921: q<=8'b00000000;
	12'h0x922: q<=8'b10101000;
	12'h0x923: q<=8'b10000100;
	12'h0x924: q<=8'b10011110;
	12'h0x925: q<=8'b10101001;
	12'h0x926: q<=8'b00001000;
	12'h0x927: q<=8'b00100000;
	12'h0x928: q<=8'b01001100;
	12'h0x929: q<=8'b11011111;
	12'h0x92a: q<=8'b10101001;
	12'h0x92b: q<=8'b00000000;
	12'h0x92c: q<=8'b00100000;
	12'h0x92d: q<=8'b01001010;
	12'h0x92e: q<=8'b11011111;
	12'h0x92f: q<=8'b00100000;
	12'h0x930: q<=8'b01100111;
	12'h0x931: q<=8'b10111001;
	12'h0x932: q<=8'b00100000;
	12'h0x933: q<=8'b00111001;
	12'h0x934: q<=8'b11011111;
	12'h0x935: q<=8'b11000110;
	12'h0x936: q<=8'b00110111;
	12'h0x937: q<=8'b00010000;
	12'h0x938: q<=8'b10101100;
	12'h0x939: q<=8'b00100000;
	12'h0x93a: q<=8'b01000100;
	12'h0x93b: q<=8'b10111001;
	12'h0x93c: q<=8'b10101001;
	12'h0x93d: q<=8'b00000001;
	12'h0x93e: q<=8'b00100000;
	12'h0x93f: q<=8'b01101010;
	12'h0x940: q<=8'b11011111;
	12'h0x941: q<=8'b00100000;
	12'h0x942: q<=8'b00001001;
	12'h0x943: q<=8'b11011111;
	12'h0x944: q<=8'b10100110;
	12'h0x945: q<=8'b01110100;
	12'h0x946: q<=8'b10100100;
	12'h0x947: q<=8'b01110101;
	12'h0x948: q<=8'b10100101;
	12'h0x949: q<=8'b01110110;
	12'h0x94a: q<=8'b10000101;
	12'h0x94b: q<=8'b01110100;
	12'h0x94c: q<=8'b10000110;
	12'h0x94d: q<=8'b01110110;
	12'h0x94e: q<=8'b10100101;
	12'h0x94f: q<=8'b01110111;
	12'h0x950: q<=8'b10000101;
	12'h0x951: q<=8'b01110101;
	12'h0x952: q<=8'b10000100;
	12'h0x953: q<=8'b01110111;
	12'h0x954: q<=8'b01100000;
	12'h0x955: q<=8'b10100101;
	12'h0x956: q<=8'b01010111;
	12'h0x957: q<=8'b01001010;
	12'h0x958: q<=8'b01001010;
	12'h0x959: q<=8'b01001010;
	12'h0x95a: q<=8'b01001010;
	12'h0x95b: q<=8'b10100000;
	12'h0x95c: q<=8'b00000000;
	12'h0x95d: q<=8'b11001000;
	12'h0x95e: q<=8'b01001010;
	12'h0x95f: q<=8'b11010000;
	12'h0x960: q<=8'b11111100;
	12'h0x961: q<=8'b00011000;
	12'h0x962: q<=8'b01101001;
	12'h0x963: q<=8'b00000010;
	12'h0x964: q<=8'b10100000;
	12'h0x965: q<=8'b00000000;
	12'h0x966: q<=8'b01100000;
	12'h0x967: q<=8'b10101101;
	12'h0x968: q<=8'b00010101;
	12'h0x969: q<=8'b00000100;
	12'h0x96a: q<=8'b11110000;
	12'h0x96b: q<=8'b00001001;
	12'h0x96c: q<=8'b10101101;
	12'h0x96d: q<=8'b01101111;
	12'h0x96e: q<=8'b11001110;
	12'h0x96f: q<=8'b10101110;
	12'h0x970: q<=8'b01101110;
	12'h0x971: q<=8'b11001110;
	12'h0x972: q<=8'b10111000;
	12'h0x973: q<=8'b01010000;
	12'h0x974: q<=8'b00000110;
	12'h0x975: q<=8'b10101101;
	12'h0x976: q<=8'b10000111;
	12'h0x977: q<=8'b11001110;
	12'h0x978: q<=8'b10101110;
	12'h0x979: q<=8'b10000110;
	12'h0x97a: q<=8'b11001110;
	12'h0x97b: q<=8'b01100000;
	12'h0x97c: q<=8'b11110000;
	12'h0x97d: q<=8'b11100111;
	12'h0x97e: q<=8'b11001111;
	12'h0x97f: q<=8'b10101010;
	12'h0x980: q<=8'b10000000;
	12'h0x981: q<=8'b01010110;
	12'h0x982: q<=8'b00110001;
	12'h0x983: q<=8'b00011001;
	12'h0x984: q<=8'b00010000;
	12'h0x985: q<=8'b00011001;
	12'h0x986: q<=8'b00110001;
	12'h0x987: q<=8'b01010110;
	12'h0x988: q<=8'b10000000;
	12'h0x989: q<=8'b10101010;
	12'h0x98a: q<=8'b11001111;
	12'h0x98b: q<=8'b11100111;
	12'h0x98c: q<=8'b11110000;
	12'h0x98d: q<=8'b11110000;
	12'h0x98e: q<=8'b11110000;
	12'h0x98f: q<=8'b10111000;
	12'h0x990: q<=8'b10000000;
	12'h0x991: q<=8'b01001000;
	12'h0x992: q<=8'b00010000;
	12'h0x993: q<=8'b00010000;
	12'h0x994: q<=8'b00010000;
	12'h0x995: q<=8'b00010000;
	12'h0x996: q<=8'b00010000;
	12'h0x997: q<=8'b01001000;
	12'h0x998: q<=8'b10000000;
	12'h0x999: q<=8'b10111000;
	12'h0x99a: q<=8'b11110000;
	12'h0x99b: q<=8'b11110000;
	12'h0x99c: q<=8'b11110000;
	12'h0x99d: q<=8'b11110000;
	12'h0x99e: q<=8'b10111000;
	12'h0x99f: q<=8'b10111000;
	12'h0x9a0: q<=8'b10000000;
	12'h0x9a1: q<=8'b01001000;
	12'h0x9a2: q<=8'b01001000;
	12'h0x9a3: q<=8'b00010000;
	12'h0x9a4: q<=8'b00010000;
	12'h0x9a5: q<=8'b00010000;
	12'h0x9a6: q<=8'b01001000;
	12'h0x9a7: q<=8'b01001000;
	12'h0x9a8: q<=8'b10000000;
	12'h0x9a9: q<=8'b10111000;
	12'h0x9aa: q<=8'b10111000;
	12'h0x9ab: q<=8'b11110000;
	12'h0x9ac: q<=8'b11101100;
	12'h0x9ad: q<=8'b11010101;
	12'h0x9ae: q<=8'b10110001;
	12'h0x9af: q<=8'b10010000;
	12'h0x9b0: q<=8'b01110000;
	12'h0x9b1: q<=8'b01001111;
	12'h0x9b2: q<=8'b00101011;
	12'h0x9b3: q<=8'b00010100;
	12'h0x9b4: q<=8'b00010100;
	12'h0x9b5: q<=8'b00101011;
	12'h0x9b6: q<=8'b01001111;
	12'h0x9b7: q<=8'b01110000;
	12'h0x9b8: q<=8'b10010000;
	12'h0x9b9: q<=8'b10110001;
	12'h0x9ba: q<=8'b11010101;
	12'h0x9bb: q<=8'b11101100;
	12'h0x9bc: q<=8'b11110000;
	12'h0x9bd: q<=8'b11000000;
	12'h0x9be: q<=8'b10100000;
	12'h0x9bf: q<=8'b10010100;
	12'h0x9c0: q<=8'b01101100;
	12'h0x9c1: q<=8'b01100000;
	12'h0x9c2: q<=8'b01000000;
	12'h0x9c3: q<=8'b00010000;
	12'h0x9c4: q<=8'b00010000;
	12'h0x9c5: q<=8'b01000000;
	12'h0x9c6: q<=8'b01100000;
	12'h0x9c7: q<=8'b01101100;
	12'h0x9c8: q<=8'b10010100;
	12'h0x9c9: q<=8'b10100000;
	12'h0x9ca: q<=8'b11000000;
	12'h0x9cb: q<=8'b11110000;
	12'h0x9cc: q<=8'b11011001;
	12'h0x9cd: q<=8'b11000010;
	12'h0x9ce: q<=8'b10101100;
	12'h0x9cf: q<=8'b10010111;
	12'h0x9d0: q<=8'b10000000;
	12'h0x9d1: q<=8'b01101001;
	12'h0x9d2: q<=8'b01010010;
	12'h0x9d3: q<=8'b00111100;
	12'h0x9d4: q<=8'b00100111;
	12'h0x9d5: q<=8'b00010000;
	12'h0x9d6: q<=8'b00110101;
	12'h0x9d7: q<=8'b01011010;
	12'h0x9d8: q<=8'b10000000;
	12'h0x9d9: q<=8'b10100110;
	12'h0x9da: q<=8'b11001010;
	12'h0x9db: q<=8'b11110000;
	12'h0x9dc: q<=8'b11101010;
	12'h0x9dd: q<=8'b11100000;
	12'h0x9de: q<=8'b10011100;
	12'h0x9df: q<=8'b10000000;
	12'h0x9e0: q<=8'b01100100;
	12'h0x9e1: q<=8'b00100000;
	12'h0x9e2: q<=8'b00010110;
	12'h0x9e3: q<=8'b01010000;
	12'h0x9e4: q<=8'b00010110;
	12'h0x9e5: q<=8'b00100000;
	12'h0x9e6: q<=8'b01100100;
	12'h0x9e7: q<=8'b10000000;
	12'h0x9e8: q<=8'b10011100;
	12'h0x9e9: q<=8'b11100000;
	12'h0x9ea: q<=8'b11101010;
	12'h0x9eb: q<=8'b10110000;
	12'h0x9ec: q<=8'b00010000;
	12'h0x9ed: q<=8'b00011110;
	12'h0x9ee: q<=8'b00101100;
	12'h0x9ef: q<=8'b00111010;
	12'h0x9f0: q<=8'b01001000;
	12'h0x9f1: q<=8'b01010110;
	12'h0x9f2: q<=8'b01100100;
	12'h0x9f3: q<=8'b01110000;
	12'h0x9f4: q<=8'b10010000;
	12'h0x9f5: q<=8'b10011110;
	12'h0x9f6: q<=8'b10101100;
	12'h0x9f7: q<=8'b10111010;
	12'h0x9f8: q<=8'b11001000;
	12'h0x9f9: q<=8'b11010110;
	12'h0x9fa: q<=8'b11100100;
	12'h0x9fb: q<=8'b11110000;
	12'h0x9fc: q<=8'b00010000;
	12'h0x9fd: q<=8'b00011110;
	12'h0x9fe: q<=8'b00101101;
	12'h0x9ff: q<=8'b00111100;
	12'h0xa00: q<=8'b01001011;
	12'h0xa01: q<=8'b01011010;
	12'h0xa02: q<=8'b01101001;
	12'h0xa03: q<=8'b01111000;
	12'h0xa04: q<=8'b10000111;
	12'h0xa05: q<=8'b10010110;
	12'h0xa06: q<=8'b10100101;
	12'h0xa07: q<=8'b10110100;
	12'h0xa08: q<=8'b11000011;
	12'h0xa09: q<=8'b11010010;
	12'h0xa0a: q<=8'b11100001;
	12'h0xa0b: q<=8'b11110000;
	12'h0xa0c: q<=8'b00010000;
	12'h0xa0d: q<=8'b00010000;
	12'h0xa0e: q<=8'b00010000;
	12'h0xa0f: q<=8'b00010000;
	12'h0xa10: q<=8'b00010110;
	12'h0xa11: q<=8'b00101001;
	12'h0xa12: q<=8'b01000110;
	12'h0xa13: q<=8'b01101001;
	12'h0xa14: q<=8'b10010111;
	12'h0xa15: q<=8'b10111010;
	12'h0xa16: q<=8'b11010111;
	12'h0xa17: q<=8'b11101010;
	12'h0xa18: q<=8'b11110000;
	12'h0xa19: q<=8'b11110000;
	12'h0xa1a: q<=8'b11110000;
	12'h0xa1b: q<=8'b11110000;
	12'h0xa1c: q<=8'b00010000;
	12'h0xa1d: q<=8'b00100100;
	12'h0xa1e: q<=8'b00110000;
	12'h0xa1f: q<=8'b00110110;
	12'h0xa20: q<=8'b00111110;
	12'h0xa21: q<=8'b01001001;
	12'h0xa22: q<=8'b01011010;
	12'h0xa23: q<=8'b01110101;
	12'h0xa24: q<=8'b10010100;
	12'h0xa25: q<=8'b10100100;
	12'h0xa26: q<=8'b10101100;
	12'h0xa27: q<=8'b10111010;
	12'h0xa28: q<=8'b11011010;
	12'h0xa29: q<=8'b11100010;
	12'h0xa2a: q<=8'b11101010;
	12'h0xa2b: q<=8'b11110000;
	12'h0xa2c: q<=8'b10000000;
	12'h0xa2d: q<=8'b01110000;
	12'h0xa2e: q<=8'b01001000;
	12'h0xa2f: q<=8'b00100000;
	12'h0xa30: q<=8'b00010000;
	12'h0xa31: q<=8'b00100000;
	12'h0xa32: q<=8'b01001000;
	12'h0xa33: q<=8'b01110000;
	12'h0xa34: q<=8'b10000000;
	12'h0xa35: q<=8'b10010000;
	12'h0xa36: q<=8'b10111000;
	12'h0xa37: q<=8'b11100000;
	12'h0xa38: q<=8'b11110000;
	12'h0xa39: q<=8'b11100000;
	12'h0xa3a: q<=8'b10111000;
	12'h0xa3b: q<=8'b10010000;
	12'h0xa3c: q<=8'b11011010;
	12'h0xa3d: q<=8'b10100100;
	12'h0xa3e: q<=8'b10000111;
	12'h0xa3f: q<=8'b10000000;
	12'h0xa40: q<=8'b01111001;
	12'h0xa41: q<=8'b01011100;
	12'h0xa42: q<=8'b00100110;
	12'h0xa43: q<=8'b00010000;
	12'h0xa44: q<=8'b00010000;
	12'h0xa45: q<=8'b00100000;
	12'h0xa46: q<=8'b01001000;
	12'h0xa47: q<=8'b10000000;
	12'h0xa48: q<=8'b10111000;
	12'h0xa49: q<=8'b11100000;
	12'h0xa4a: q<=8'b11110000;
	12'h0xa4b: q<=8'b11110000;
	12'h0xa4c: q<=8'b00010000;
	12'h0xa4d: q<=8'b00010000;
	12'h0xa4e: q<=8'b00110000;
	12'h0xa4f: q<=8'b00110000;
	12'h0xa50: q<=8'b01010000;
	12'h0xa51: q<=8'b01010000;
	12'h0xa52: q<=8'b01110000;
	12'h0xa53: q<=8'b01110000;
	12'h0xa54: q<=8'b10010000;
	12'h0xa55: q<=8'b10010000;
	12'h0xa56: q<=8'b10110000;
	12'h0xa57: q<=8'b10110000;
	12'h0xa58: q<=8'b11010000;
	12'h0xa59: q<=8'b11010000;
	12'h0xa5a: q<=8'b11110000;
	12'h0xa5b: q<=8'b11110000;
	12'h0xa5c: q<=8'b10110000;
	12'h0xa5d: q<=8'b10000000;
	12'h0xa5e: q<=8'b01010000;
	12'h0xa5f: q<=8'b01000111;
	12'h0xa60: q<=8'b00011000;
	12'h0xa61: q<=8'b00110000;
	12'h0xa62: q<=8'b00011000;
	12'h0xa63: q<=8'b01000111;
	12'h0xa64: q<=8'b01010000;
	12'h0xa65: q<=8'b10000000;
	12'h0xa66: q<=8'b10110000;
	12'h0xa67: q<=8'b10111001;
	12'h0xa68: q<=8'b11101000;
	12'h0xa69: q<=8'b11010100;
	12'h0xa6a: q<=8'b11101000;
	12'h0xa6b: q<=8'b10111001;
	12'h0xa6c: q<=8'b00010000;
	12'h0xa6d: q<=8'b00011110;
	12'h0xa6e: q<=8'b00100001;
	12'h0xa6f: q<=8'b00101000;
	12'h0xa70: q<=8'b00111100;
	12'h0xa71: q<=8'b01010101;
	12'h0xa72: q<=8'b01100110;
	12'h0xa73: q<=8'b01110011;
	12'h0xa74: q<=8'b10001101;
	12'h0xa75: q<=8'b10011010;
	12'h0xa76: q<=8'b10101011;
	12'h0xa77: q<=8'b11000100;
	12'h0xa78: q<=8'b11011000;
	12'h0xa79: q<=8'b11011111;
	12'h0xa7a: q<=8'b11100010;
	12'h0xa7b: q<=8'b11110000;
	12'h0xa7c: q<=8'b10000000;
	12'h0xa7d: q<=8'b10101010;
	12'h0xa7e: q<=8'b11001111;
	12'h0xa7f: q<=8'b11100111;
	12'h0xa80: q<=8'b11110000;
	12'h0xa81: q<=8'b11100111;
	12'h0xa82: q<=8'b11001111;
	12'h0xa83: q<=8'b10101010;
	12'h0xa84: q<=8'b10000000;
	12'h0xa85: q<=8'b01010110;
	12'h0xa86: q<=8'b00110001;
	12'h0xa87: q<=8'b00011001;
	12'h0xa88: q<=8'b00010000;
	12'h0xa89: q<=8'b00011001;
	12'h0xa8a: q<=8'b00110001;
	12'h0xa8b: q<=8'b01010110;
	12'h0xa8c: q<=8'b10000000;
	12'h0xa8d: q<=8'b10111000;
	12'h0xa8e: q<=8'b11110000;
	12'h0xa8f: q<=8'b11110000;
	12'h0xa90: q<=8'b11110000;
	12'h0xa91: q<=8'b11110000;
	12'h0xa92: q<=8'b11110000;
	12'h0xa93: q<=8'b10111000;
	12'h0xa94: q<=8'b10000000;
	12'h0xa95: q<=8'b01001000;
	12'h0xa96: q<=8'b00010000;
	12'h0xa97: q<=8'b00010000;
	12'h0xa98: q<=8'b00010000;
	12'h0xa99: q<=8'b00010000;
	12'h0xa9a: q<=8'b00010000;
	12'h0xa9b: q<=8'b01001000;
	12'h0xa9c: q<=8'b10000000;
	12'h0xa9d: q<=8'b10111000;
	12'h0xa9e: q<=8'b10111000;
	12'h0xa9f: q<=8'b11110000;
	12'h0xaa0: q<=8'b11110000;
	12'h0xaa1: q<=8'b11110000;
	12'h0xaa2: q<=8'b10111000;
	12'h0xaa3: q<=8'b10111000;
	12'h0xaa4: q<=8'b10000000;
	12'h0xaa5: q<=8'b01001000;
	12'h0xaa6: q<=8'b01001000;
	12'h0xaa7: q<=8'b00010000;
	12'h0xaa8: q<=8'b00010000;
	12'h0xaa9: q<=8'b00010000;
	12'h0xaaa: q<=8'b01001000;
	12'h0xaab: q<=8'b01001000;
	12'h0xaac: q<=8'b10010100;
	12'h0xaad: q<=8'b10110000;
	12'h0xaae: q<=8'b10111000;
	12'h0xaaf: q<=8'b10100111;
	12'h0xab0: q<=8'b10100111;
	12'h0xab1: q<=8'b10111000;
	12'h0xab2: q<=8'b10110000;
	12'h0xab3: q<=8'b10010100;
	12'h0xab4: q<=8'b01101100;
	12'h0xab5: q<=8'b01010000;
	12'h0xab6: q<=8'b01001000;
	12'h0xab7: q<=8'b01011001;
	12'h0xab8: q<=8'b01011001;
	12'h0xab9: q<=8'b01001000;
	12'h0xaba: q<=8'b01010000;
	12'h0xabb: q<=8'b01101100;
	12'h0xabc: q<=8'b10010110;
	12'h0xabd: q<=8'b10100011;
	12'h0xabe: q<=8'b11000101;
	12'h0xabf: q<=8'b11110000;
	12'h0xac0: q<=8'b11110000;
	12'h0xac1: q<=8'b11000101;
	12'h0xac2: q<=8'b10100011;
	12'h0xac3: q<=8'b10010110;
	12'h0xac4: q<=8'b01101010;
	12'h0xac5: q<=8'b01011101;
	12'h0xac6: q<=8'b00111011;
	12'h0xac7: q<=8'b00010000;
	12'h0xac8: q<=8'b00010000;
	12'h0xac9: q<=8'b00111011;
	12'h0xaca: q<=8'b01011101;
	12'h0xacb: q<=8'b01101010;
	12'h0xacc: q<=8'b00111101;
	12'h0xacd: q<=8'b01101010;
	12'h0xace: q<=8'b10010111;
	12'h0xacf: q<=8'b11000100;
	12'h0xad0: q<=8'b11110000;
	12'h0xad1: q<=8'b11000100;
	12'h0xad2: q<=8'b10010111;
	12'h0xad3: q<=8'b01101010;
	12'h0xad4: q<=8'b00111101;
	12'h0xad5: q<=8'b00010000;
	12'h0xad6: q<=8'b00010000;
	12'h0xad7: q<=8'b00010000;
	12'h0xad8: q<=8'b00010000;
	12'h0xad9: q<=8'b00010000;
	12'h0xada: q<=8'b00010000;
	12'h0xadb: q<=8'b00010000;
	12'h0xadc: q<=8'b10100000;
	12'h0xadd: q<=8'b11100000;
	12'h0xade: q<=8'b11101010;
	12'h0xadf: q<=8'b10110000;
	12'h0xae0: q<=8'b11101010;
	12'h0xae1: q<=8'b11100000;
	12'h0xae2: q<=8'b10100000;
	12'h0xae3: q<=8'b10000000;
	12'h0xae4: q<=8'b01100000;
	12'h0xae5: q<=8'b00100000;
	12'h0xae6: q<=8'b00010110;
	12'h0xae7: q<=8'b01010000;
	12'h0xae8: q<=8'b00010110;
	12'h0xae9: q<=8'b00100000;
	12'h0xaea: q<=8'b01100000;
	12'h0xaeb: q<=8'b10000000;
	12'h0xaec: q<=8'b11110000;
	12'h0xaed: q<=8'b11010000;
	12'h0xaee: q<=8'b10110000;
	12'h0xaef: q<=8'b10010000;
	12'h0xaf0: q<=8'b01110000;
	12'h0xaf1: q<=8'b01010000;
	12'h0xaf2: q<=8'b00110000;
	12'h0xaf3: q<=8'b00010000;
	12'h0xaf4: q<=8'b00010000;
	12'h0xaf5: q<=8'b00110000;
	12'h0xaf6: q<=8'b01010000;
	12'h0xaf7: q<=8'b01110000;
	12'h0xaf8: q<=8'b10010000;
	12'h0xaf9: q<=8'b10110000;
	12'h0xafa: q<=8'b11010000;
	12'h0xafb: q<=8'b11110000;
	12'h0xafc: q<=8'b01000000;
	12'h0xafd: q<=8'b01000000;
	12'h0xafe: q<=8'b01000000;
	12'h0xaff: q<=8'b01000000;
	12'h0xb00: q<=8'b01000000;
	12'h0xb01: q<=8'b01000000;
	12'h0xb02: q<=8'b01000000;
	12'h0xb03: q<=8'b01000000;
	12'h0xb04: q<=8'b01000000;
	12'h0xb05: q<=8'b01000000;
	12'h0xb06: q<=8'b01000000;
	12'h0xb07: q<=8'b01000000;
	12'h0xb08: q<=8'b01000000;
	12'h0xb09: q<=8'b01000000;
	12'h0xb0a: q<=8'b01000000;
	12'h0xb0b: q<=8'b01000000;
	12'h0xb0c: q<=8'b11110000;
	12'h0xb0d: q<=8'b11001011;
	12'h0xb0e: q<=8'b10100110;
	12'h0xb0f: q<=8'b10000000;
	12'h0xb10: q<=8'b01011100;
	12'h0xb11: q<=8'b00111001;
	12'h0xb12: q<=8'b00100000;
	12'h0xb13: q<=8'b00010010;
	12'h0xb14: q<=8'b00010010;
	12'h0xb15: q<=8'b00100000;
	12'h0xb16: q<=8'b00111001;
	12'h0xb17: q<=8'b01011100;
	12'h0xb18: q<=8'b10000000;
	12'h0xb19: q<=8'b10100110;
	12'h0xb1a: q<=8'b11001011;
	12'h0xb1b: q<=8'b11110000;
	12'h0xb1c: q<=8'b11000000;
	12'h0xb1d: q<=8'b10100110;
	12'h0xb1e: q<=8'b10001010;
	12'h0xb1f: q<=8'b01101010;
	12'h0xb20: q<=8'b01001010;
	12'h0xb21: q<=8'b00101111;
	12'h0xb22: q<=8'b00010100;
	12'h0xb23: q<=8'b00100100;
	12'h0xb24: q<=8'b00100000;
	12'h0xb25: q<=8'b00111001;
	12'h0xb26: q<=8'b01011001;
	12'h0xb27: q<=8'b01110101;
	12'h0xb28: q<=8'b01110010;
	12'h0xb29: q<=8'b10010000;
	12'h0xb2a: q<=8'b10110000;
	12'h0xb2b: q<=8'b11010000;
	12'h0xb2c: q<=8'b10000000;
	12'h0xb2d: q<=8'b01010111;
	12'h0xb2e: q<=8'b01001000;
	12'h0xb2f: q<=8'b01010111;
	12'h0xb30: q<=8'b10000000;
	12'h0xb31: q<=8'b10101001;
	12'h0xb32: q<=8'b10111010;
	12'h0xb33: q<=8'b10101001;
	12'h0xb34: q<=8'b10000000;
	12'h0xb35: q<=8'b01010111;
	12'h0xb36: q<=8'b01001000;
	12'h0xb37: q<=8'b01010111;
	12'h0xb38: q<=8'b10000000;
	12'h0xb39: q<=8'b10101001;
	12'h0xb3a: q<=8'b10111010;
	12'h0xb3b: q<=8'b10101001;
	12'h0xb3c: q<=8'b11100100;
	12'h0xb3d: q<=8'b11101000;
	12'h0xb3e: q<=8'b10110111;
	12'h0xb3f: q<=8'b10000000;
	12'h0xb40: q<=8'b10110111;
	12'h0xb41: q<=8'b11101000;
	12'h0xb42: q<=8'b11100100;
	12'h0xb43: q<=8'b10110010;
	12'h0xb44: q<=8'b01111010;
	12'h0xb45: q<=8'b01000111;
	12'h0xb46: q<=8'b00100000;
	12'h0xb47: q<=8'b00010000;
	12'h0xb48: q<=8'b00100000;
	12'h0xb49: q<=8'b01000111;
	12'h0xb4a: q<=8'b01111010;
	12'h0xb4b: q<=8'b10110010;
	12'h0xb4c: q<=8'b10010000;
	12'h0xb4d: q<=8'b01110000;
	12'h0xb4e: q<=8'b01110000;
	12'h0xb4f: q<=8'b01010000;
	12'h0xb50: q<=8'b01010000;
	12'h0xb51: q<=8'b00110000;
	12'h0xb52: q<=8'b00110000;
	12'h0xb53: q<=8'b00010000;
	12'h0xb54: q<=8'b00010000;
	12'h0xb55: q<=8'b00110000;
	12'h0xb56: q<=8'b00110000;
	12'h0xb57: q<=8'b01010000;
	12'h0xb58: q<=8'b01010000;
	12'h0xb59: q<=8'b01110000;
	12'h0xb5a: q<=8'b01110000;
	12'h0xb5b: q<=8'b10010000;
	12'h0xb5c: q<=8'b11100110;
	12'h0xb5d: q<=8'b11010000;
	12'h0xb5e: q<=8'b11100110;
	12'h0xb5f: q<=8'b10111001;
	12'h0xb60: q<=8'b10101110;
	12'h0xb61: q<=8'b10000000;
	12'h0xb62: q<=8'b01010010;
	12'h0xb63: q<=8'b01000111;
	12'h0xb64: q<=8'b00010100;
	12'h0xb65: q<=8'b00110000;
	12'h0xb66: q<=8'b00010100;
	12'h0xb67: q<=8'b01000111;
	12'h0xb68: q<=8'b01010010;
	12'h0xb69: q<=8'b10000000;
	12'h0xb6a: q<=8'b10101110;
	12'h0xb6b: q<=8'b10111001;
	12'h0xb6c: q<=8'b01111110;
	12'h0xb6d: q<=8'b01101010;
	12'h0xb6e: q<=8'b01010001;
	12'h0xb6f: q<=8'b00111010;
	12'h0xb70: q<=8'b00101100;
	12'h0xb71: q<=8'b00101100;
	12'h0xb72: q<=8'b00111000;
	12'h0xb73: q<=8'b01001110;
	12'h0xb74: q<=8'b01001110;
	12'h0xb75: q<=8'b00111000;
	12'h0xb76: q<=8'b00101100;
	12'h0xb77: q<=8'b00101100;
	12'h0xb78: q<=8'b00111010;
	12'h0xb79: q<=8'b01010001;
	12'h0xb7a: q<=8'b01101010;
	12'h0xb7b: q<=8'b01111110;
	12'h0xb7c: q<=8'b00000101;
	12'h0xb7d: q<=8'b00000110;
	12'h0xb7e: q<=8'b00000111;
	12'h0xb7f: q<=8'b00001000;
	12'h0xb80: q<=8'b00001001;
	12'h0xb81: q<=8'b00001010;
	12'h0xb82: q<=8'b00001011;
	12'h0xb83: q<=8'b00001100;
	12'h0xb84: q<=8'b00001101;
	12'h0xb85: q<=8'b00001110;
	12'h0xb86: q<=8'b00001111;
	12'h0xb87: q<=8'b00000000;
	12'h0xb88: q<=8'b00000001;
	12'h0xb89: q<=8'b00000010;
	12'h0xb8a: q<=8'b00000011;
	12'h0xb8b: q<=8'b00000100;
	12'h0xb8c: q<=8'b00000100;
	12'h0xb8d: q<=8'b00000100;
	12'h0xb8e: q<=8'b00001000;
	12'h0xb8f: q<=8'b00001000;
	12'h0xb90: q<=8'b00001000;
	12'h0xb91: q<=8'b00001000;
	12'h0xb92: q<=8'b00001100;
	12'h0xb93: q<=8'b00001100;
	12'h0xb94: q<=8'b00001100;
	12'h0xb95: q<=8'b00001100;
	12'h0xb96: q<=8'b00000000;
	12'h0xb97: q<=8'b00000000;
	12'h0xb98: q<=8'b00000000;
	12'h0xb99: q<=8'b00000000;
	12'h0xb9a: q<=8'b00000100;
	12'h0xb9b: q<=8'b00000100;
	12'h0xb9c: q<=8'b00000100;
	12'h0xb9d: q<=8'b00001000;
	12'h0xb9e: q<=8'b00000100;
	12'h0xb9f: q<=8'b00001000;
	12'h0xba0: q<=8'b00001000;
	12'h0xba1: q<=8'b00001100;
	12'h0xba2: q<=8'b00001000;
	12'h0xba3: q<=8'b00001100;
	12'h0xba4: q<=8'b00001100;
	12'h0xba5: q<=8'b00000000;
	12'h0xba6: q<=8'b00001100;
	12'h0xba7: q<=8'b00000000;
	12'h0xba8: q<=8'b00000000;
	12'h0xba9: q<=8'b00000100;
	12'h0xbaa: q<=8'b00000000;
	12'h0xbab: q<=8'b00000100;
	12'h0xbac: q<=8'b00000110;
	12'h0xbad: q<=8'b00000111;
	12'h0xbae: q<=8'b00001001;
	12'h0xbaf: q<=8'b00001000;
	12'h0xbb0: q<=8'b00000111;
	12'h0xbb1: q<=8'b00001001;
	12'h0xbb2: q<=8'b00001010;
	12'h0xbb3: q<=8'b00001100;
	12'h0xbb4: q<=8'b00001110;
	12'h0xbb5: q<=8'b00001111;
	12'h0xbb6: q<=8'b00000001;
	12'h0xbb7: q<=8'b00000000;
	12'h0xbb8: q<=8'b00001111;
	12'h0xbb9: q<=8'b00000001;
	12'h0xbba: q<=8'b00000010;
	12'h0xbbb: q<=8'b00000100;
	12'h0xbbc: q<=8'b00000111;
	12'h0xbbd: q<=8'b00000110;
	12'h0xbbe: q<=8'b00000101;
	12'h0xbbf: q<=8'b00001000;
	12'h0xbc0: q<=8'b00001011;
	12'h0xbc1: q<=8'b00001010;
	12'h0xbc2: q<=8'b00001001;
	12'h0xbc3: q<=8'b00001100;
	12'h0xbc4: q<=8'b00001111;
	12'h0xbc5: q<=8'b00001110;
	12'h0xbc6: q<=8'b00001101;
	12'h0xbc7: q<=8'b00000000;
	12'h0xbc8: q<=8'b00000011;
	12'h0xbc9: q<=8'b00000010;
	12'h0xbca: q<=8'b00000001;
	12'h0xbcb: q<=8'b00000100;
	12'h0xbcc: q<=8'b00000101;
	12'h0xbcd: q<=8'b00000101;
	12'h0xbce: q<=8'b00000101;
	12'h0xbcf: q<=8'b00000101;
	12'h0xbd0: q<=8'b00001011;
	12'h0xbd1: q<=8'b00001011;
	12'h0xbd2: q<=8'b00001011;
	12'h0xbd3: q<=8'b00001011;
	12'h0xbd4: q<=8'b00001011;
	12'h0xbd5: q<=8'b00000000;
	12'h0xbd6: q<=8'b00000000;
	12'h0xbd7: q<=8'b00000000;
	12'h0xbd8: q<=8'b00000000;
	12'h0xbd9: q<=8'b00000000;
	12'h0xbda: q<=8'b00000000;
	12'h0xbdb: q<=8'b00000101;
	12'h0xbdc: q<=8'b00000100;
	12'h0xbdd: q<=8'b00001000;
	12'h0xbde: q<=8'b00001011;
	12'h0xbdf: q<=8'b00000101;
	12'h0xbe0: q<=8'b00001000;
	12'h0xbe1: q<=8'b00001100;
	12'h0xbe2: q<=8'b00001110;
	12'h0xbe3: q<=8'b00001001;
	12'h0xbe4: q<=8'b00001100;
	12'h0xbe5: q<=8'b00000000;
	12'h0xbe6: q<=8'b00000011;
	12'h0xbe7: q<=8'b00001101;
	12'h0xbe8: q<=8'b00000000;
	12'h0xbe9: q<=8'b00000100;
	12'h0xbea: q<=8'b00000111;
	12'h0xbeb: q<=8'b00000010;
	12'h0xbec: q<=8'b00001101;
	12'h0xbed: q<=8'b00001101;
	12'h0xbee: q<=8'b00001101;
	12'h0xbef: q<=8'b00001101;
	12'h0xbf0: q<=8'b00001101;
	12'h0xbf1: q<=8'b00001101;
	12'h0xbf2: q<=8'b00001101;
	12'h0xbf3: q<=8'b00000000;
	12'h0xbf4: q<=8'b00000011;
	12'h0xbf5: q<=8'b00000011;
	12'h0xbf6: q<=8'b00000011;
	12'h0xbf7: q<=8'b00000011;
	12'h0xbf8: q<=8'b00000011;
	12'h0xbf9: q<=8'b00000011;
	12'h0xbfa: q<=8'b00000011;
	12'h0xbfb: q<=8'b00000000;
	12'h0xbfc: q<=8'b00000000;
	12'h0xbfd: q<=8'b00000000;
	12'h0xbfe: q<=8'b00000000;
	12'h0xbff: q<=8'b00000000;
	12'h0xc00: q<=8'b00000000;
	12'h0xc01: q<=8'b00000000;
	12'h0xc02: q<=8'b00000000;
	12'h0xc03: q<=8'b00000000;
	12'h0xc04: q<=8'b00000000;
	12'h0xc05: q<=8'b00000000;
	12'h0xc06: q<=8'b00000000;
	12'h0xc07: q<=8'b00000000;
	12'h0xc08: q<=8'b00000000;
	12'h0xc09: q<=8'b00000000;
	12'h0xc0a: q<=8'b00000000;
	12'h0xc0b: q<=8'b00000000;
	12'h0xc0c: q<=8'b00001100;
	12'h0xc0d: q<=8'b00001100;
	12'h0xc0e: q<=8'b00001100;
	12'h0xc0f: q<=8'b00001101;
	12'h0xc10: q<=8'b00001110;
	12'h0xc11: q<=8'b00001111;
	12'h0xc12: q<=8'b00001111;
	12'h0xc13: q<=8'b00000000;
	12'h0xc14: q<=8'b00000001;
	12'h0xc15: q<=8'b00000001;
	12'h0xc16: q<=8'b00000010;
	12'h0xc17: q<=8'b00000011;
	12'h0xc18: q<=8'b00000100;
	12'h0xc19: q<=8'b00000100;
	12'h0xc1a: q<=8'b00000100;
	12'h0xc1b: q<=8'b00000000;
	12'h0xc1c: q<=8'b00001110;
	12'h0xc1d: q<=8'b00001101;
	12'h0xc1e: q<=8'b00001100;
	12'h0xc1f: q<=8'b00001101;
	12'h0xc20: q<=8'b00001101;
	12'h0xc21: q<=8'b00001101;
	12'h0xc22: q<=8'b00000001;
	12'h0xc23: q<=8'b00001111;
	12'h0xc24: q<=8'b00000010;
	12'h0xc25: q<=8'b00000011;
	12'h0xc26: q<=8'b00000011;
	12'h0xc27: q<=8'b00000000;
	12'h0xc28: q<=8'b00000011;
	12'h0xc29: q<=8'b00000011;
	12'h0xc2a: q<=8'b00000011;
	12'h0xc2b: q<=8'b00000000;
	12'h0xc2c: q<=8'b00001011;
	12'h0xc2d: q<=8'b00001001;
	12'h0xc2e: q<=8'b00000111;
	12'h0xc2f: q<=8'b00000101;
	12'h0xc30: q<=8'b00000011;
	12'h0xc31: q<=8'b00000001;
	12'h0xc32: q<=8'b00001111;
	12'h0xc33: q<=8'b00001101;
	12'h0xc34: q<=8'b00001101;
	12'h0xc35: q<=8'b00001111;
	12'h0xc36: q<=8'b00000001;
	12'h0xc37: q<=8'b00000011;
	12'h0xc38: q<=8'b00000101;
	12'h0xc39: q<=8'b00000111;
	12'h0xc3a: q<=8'b00001001;
	12'h0xc3b: q<=8'b00001011;
	12'h0xc3c: q<=8'b00001000;
	12'h0xc3d: q<=8'b00001011;
	12'h0xc3e: q<=8'b00001100;
	12'h0xc3f: q<=8'b00000100;
	12'h0xc40: q<=8'b00000101;
	12'h0xc41: q<=8'b00001000;
	12'h0xc42: q<=8'b00001011;
	12'h0xc43: q<=8'b00001100;
	12'h0xc44: q<=8'b00001101;
	12'h0xc45: q<=8'b00001110;
	12'h0xc46: q<=8'b00001111;
	12'h0xc47: q<=8'b00000001;
	12'h0xc48: q<=8'b00000010;
	12'h0xc49: q<=8'b00000011;
	12'h0xc4a: q<=8'b00000100;
	12'h0xc4b: q<=8'b00000101;
	12'h0xc4c: q<=8'b00001100;
	12'h0xc4d: q<=8'b00000000;
	12'h0xc4e: q<=8'b00001100;
	12'h0xc4f: q<=8'b00000000;
	12'h0xc50: q<=8'b00001100;
	12'h0xc51: q<=8'b00000000;
	12'h0xc52: q<=8'b00001100;
	12'h0xc53: q<=8'b00000000;
	12'h0xc54: q<=8'b00000100;
	12'h0xc55: q<=8'b00000000;
	12'h0xc56: q<=8'b00000100;
	12'h0xc57: q<=8'b00000000;
	12'h0xc58: q<=8'b00000100;
	12'h0xc59: q<=8'b00000000;
	12'h0xc5a: q<=8'b00000100;
	12'h0xc5b: q<=8'b00000000;
	12'h0xc5c: q<=8'b00001010;
	12'h0xc5d: q<=8'b00000110;
	12'h0xc5e: q<=8'b00001100;
	12'h0xc5f: q<=8'b00001000;
	12'h0xc60: q<=8'b00001110;
	12'h0xc61: q<=8'b00001010;
	12'h0xc62: q<=8'b00000000;
	12'h0xc63: q<=8'b00001100;
	12'h0xc64: q<=8'b00000010;
	12'h0xc65: q<=8'b00001110;
	12'h0xc66: q<=8'b00000100;
	12'h0xc67: q<=8'b00000000;
	12'h0xc68: q<=8'b00000110;
	12'h0xc69: q<=8'b00000010;
	12'h0xc6a: q<=8'b00001000;
	12'h0xc6b: q<=8'b00000100;
	12'h0xc6c: q<=8'b00001110;
	12'h0xc6d: q<=8'b00001100;
	12'h0xc6e: q<=8'b00001101;
	12'h0xc6f: q<=8'b00001110;
	12'h0xc70: q<=8'b00000000;
	12'h0xc71: q<=8'b00000010;
	12'h0xc72: q<=8'b00000010;
	12'h0xc73: q<=8'b00000000;
	12'h0xc74: q<=8'b00001110;
	12'h0xc75: q<=8'b00001110;
	12'h0xc76: q<=8'b00000000;
	12'h0xc77: q<=8'b00000010;
	12'h0xc78: q<=8'b00000011;
	12'h0xc79: q<=8'b00000100;
	12'h0xc7a: q<=8'b00000010;
	12'h0xc7b: q<=8'b00000000;
	12'h0xc7c: q<=8'b00000000;
	12'h0xc7d: q<=8'b00000001;
	12'h0xc7e: q<=8'b00000010;
	12'h0xc7f: q<=8'b00000011;
	12'h0xc80: q<=8'b00000100;
	12'h0xc81: q<=8'b00000101;
	12'h0xc82: q<=8'b00000110;
	12'h0xc83: q<=8'b00000111;
	12'h0xc84: q<=8'b00001101;
	12'h0xc85: q<=8'b00001001;
	12'h0xc86: q<=8'b00001000;
	12'h0xc87: q<=8'b00001100;
	12'h0xc88: q<=8'b00001110;
	12'h0xc89: q<=8'b00001111;
	12'h0xc8a: q<=8'b00001010;
	12'h0xc8b: q<=8'b00001011;
	12'h0xc8c: q<=8'b00011000;
	12'h0xc8d: q<=8'b00011100;
	12'h0xc8e: q<=8'b00011000;
	12'h0xc8f: q<=8'b00001111;
	12'h0xc90: q<=8'b00011000;
	12'h0xc91: q<=8'b00011000;
	12'h0xc92: q<=8'b00011000;
	12'h0xc93: q<=8'b00011000;
	12'h0xc94: q<=8'b00001010;
	12'h0xc95: q<=8'b00011000;
	12'h0xc96: q<=8'b00010000;
	12'h0xc97: q<=8'b00001111;
	12'h0xc98: q<=8'b00011000;
	12'h0xc99: q<=8'b00001100;
	12'h0xc9a: q<=8'b00010100;
	12'h0xc9b: q<=8'b00001010;
	12'h0xc9c: q<=8'b01010000;
	12'h0xc9d: q<=8'b01010000;
	12'h0xc9e: q<=8'b01010000;
	12'h0xc9f: q<=8'b01101000;
	12'h0xca0: q<=8'b01010000;
	12'h0xca1: q<=8'b01010000;
	12'h0xca2: q<=8'b01101000;
	12'h0xca3: q<=8'b10110000;
	12'h0xca4: q<=8'b10100000;
	12'h0xca5: q<=8'b01010000;
	12'h0xca6: q<=8'b10010000;
	12'h0xca7: q<=8'b10000000;
	12'h0xca8: q<=8'b00100000;
	12'h0xca9: q<=8'b10110000;
	12'h0xcaa: q<=8'b01100000;
	12'h0xcab: q<=8'b10100000;
	12'h0xcac: q<=8'b01000000;
	12'h0xcad: q<=8'b00100000;
	12'h0xcae: q<=8'b01000000;
	12'h0xcaf: q<=8'b10000000;
	12'h0xcb0: q<=8'b01000000;
	12'h0xcb1: q<=8'b01000000;
	12'h0xcb2: q<=8'b01110000;
	12'h0xcb3: q<=8'b01100000;
	12'h0xcb4: q<=8'b00000000;
	12'h0xcb5: q<=8'b00100000;
	12'h0xcb6: q<=8'b01000000;
	12'h0xcb7: q<=8'b00000000;
	12'h0xcb8: q<=8'b10100000;
	12'h0xcb9: q<=8'b01000000;
	12'h0xcba: q<=8'b01000000;
	12'h0xcbb: q<=8'b00000000;
	12'h0xcbc: q<=8'b11111111;
	12'h0xcbd: q<=8'b11111111;
	12'h0xcbe: q<=8'b11111111;
	12'h0xcbf: q<=8'b11111111;
	12'h0xcc0: q<=8'b11111111;
	12'h0xcc1: q<=8'b11111111;
	12'h0xcc2: q<=8'b11111111;
	12'h0xcc3: q<=8'b00000000;
	12'h0xcc4: q<=8'b00000001;
	12'h0xcc5: q<=8'b11111111;
	12'h0xcc6: q<=8'b00000000;
	12'h0xcc7: q<=8'b00000000;
	12'h0xcc8: q<=8'b11111110;
	12'h0xcc9: q<=8'b00000001;
	12'h0xcca: q<=8'b11111111;
	12'h0xccb: q<=8'b00000001;
	12'h0xccc: q<=8'b00000000;
	12'h0xccd: q<=8'b00000000;
	12'h0xcce: q<=8'b00000000;
	12'h0xccf: q<=8'b00000000;
	12'h0xcd0: q<=8'b00000000;
	12'h0xcd1: q<=8'b00000000;
	12'h0xcd2: q<=8'b00000000;
	12'h0xcd3: q<=8'b11111111;
	12'h0xcd4: q<=8'b11111111;
	12'h0xcd5: q<=8'b11111111;
	12'h0xcd6: q<=8'b11111111;
	12'h0xcd7: q<=8'b00000000;
	12'h0xcd8: q<=8'b00000000;
	12'h0xcd9: q<=8'b11111111;
	12'h0xcda: q<=8'b00000000;
	12'h0xcdb: q<=8'b11111111;
	12'h0xcdc: q<=8'b00000000;
	12'h0xcdd: q<=8'b00000000;
	12'h0xcde: q<=8'b01100000;
	12'h0xcdf: q<=8'b01000000;
	12'h0xce0: q<=8'b00000000;
	12'h0xce1: q<=8'b00000000;
	12'h0xce2: q<=8'b01001000;
	12'h0xce3: q<=8'b01000000;
	12'h0xce4: q<=8'b01010000;
	12'h0xce5: q<=8'b00101000;
	12'h0xce6: q<=8'b01010000;
	12'h0xce7: q<=8'b00000000;
	12'h0xce8: q<=8'b00000000;
	12'h0xce9: q<=8'b01010000;
	12'h0xcea: q<=8'b00000000;
	12'h0xceb: q<=8'b01000000;
	12'h0xcec: q<=8'b00000100;
	12'h0xced: q<=8'b00000100;
	12'h0xcee: q<=8'b00000011;
	12'h0xcef: q<=8'b00000100;
	12'h0xcf0: q<=8'b00000100;
	12'h0xcf1: q<=8'b00000100;
	12'h0xcf2: q<=8'b00000011;
	12'h0xcf3: q<=8'b00000100;
	12'h0xcf4: q<=8'b00000101;
	12'h0xcf5: q<=8'b00000100;
	12'h0xcf6: q<=8'b00000100;
	12'h0xcf7: q<=8'b00000100;
	12'h0xcf8: q<=8'b00000100;
	12'h0xcf9: q<=8'b00000100;
	12'h0xcfa: q<=8'b00000100;
	12'h0xcfb: q<=8'b00000101;
	12'h0xcfc: q<=8'b00111110;
	12'h0xcfd: q<=8'b10000101;
	12'h0xcfe: q<=8'b01010101;
	12'h0xcff: q<=8'b10111001;
	12'h0xd00: q<=8'b00110101;
	12'h0xd01: q<=8'b00000100;
	12'h0xd02: q<=8'b10000101;
	12'h0xd03: q<=8'b01010110;
	12'h0xd04: q<=8'b10111001;
	12'h0xd05: q<=8'b01000101;
	12'h0xd06: q<=8'b00000100;
	12'h0xd07: q<=8'b10000101;
	12'h0xd08: q<=8'b01011000;
	12'h0xd09: q<=8'b00100000;
	12'h0xd0a: q<=8'b10011000;
	12'h0xd0b: q<=8'b11000000;
	12'h0xd0c: q<=8'b10100010;
	12'h0xd0d: q<=8'b01100001;
	12'h0xd0e: q<=8'b00100000;
	12'h0xd0f: q<=8'b01100101;
	12'h0xd10: q<=8'b11000111;
	12'h0xd11: q<=8'b10101001;
	12'h0xd12: q<=8'b00000000;
	12'h0xd13: q<=8'b10000101;
	12'h0xd14: q<=8'b10101001;
	12'h0xd15: q<=8'b00100000;
	12'h0xd16: q<=8'b00111110;
	12'h0xd17: q<=8'b10111101;
	12'h0xd18: q<=8'b10100101;
	12'h0xd19: q<=8'b01111000;
	12'h0xd1a: q<=8'b01001001;
	12'h0xd1b: q<=8'b00000111;
	12'h0xd1c: q<=8'b00001010;
	12'h0xd1d: q<=8'b11001001;
	12'h0xd1e: q<=8'b00001010;
	12'h0xd1f: q<=8'b10110000;
	12'h0xd20: q<=8'b00000010;
	12'h0xd21: q<=8'b10101001;
	12'h0xd22: q<=8'b00001010;
	12'h0xd23: q<=8'b00001010;
	12'h0xd24: q<=8'b00001010;
	12'h0xd25: q<=8'b00001010;
	12'h0xd26: q<=8'b00001010;
	12'h0xd27: q<=8'b10010001;
	12'h0xd28: q<=8'b01110100;
	12'h0xd29: q<=8'b11001000;
	12'h0xd2a: q<=8'b10101001;
	12'h0xd2b: q<=8'b01100000;
	12'h0xd2c: q<=8'b10010001;
	12'h0xd2d: q<=8'b01110100;
	12'h0xd2e: q<=8'b11001000;
	12'h0xd2f: q<=8'b10000100;
	12'h0xd30: q<=8'b10101001;
	12'h0xd31: q<=8'b10100100;
	12'h0xd32: q<=8'b01010101;
	12'h0xd33: q<=8'b10111110;
	12'h0xd34: q<=8'b11001001;
	12'h0xd35: q<=8'b11001110;
	12'h0xd36: q<=8'b10111001;
	12'h0xd37: q<=8'b11001000;
	12'h0xd38: q<=8'b11001110;
	12'h0xd39: q<=8'b10100100;
	12'h0xd3a: q<=8'b10101001;
	12'h0xd3b: q<=8'b01001100;
	12'h0xd3c: q<=8'b01011001;
	12'h0xd3d: q<=8'b11011111;
	12'h0xd3e: q<=8'b10100101;
	12'h0xd3f: q<=8'b01010111;
	12'h0xd40: q<=8'b11001001;
	12'h0xd41: q<=8'b00010000;
	12'h0xd42: q<=8'b10010000;
	12'h0xd43: q<=8'b01001000;
	12'h0xd44: q<=8'b00111000;
	12'h0xd45: q<=8'b11100101;
	12'h0xd46: q<=8'b01011111;
	12'h0xd47: q<=8'b10001101;
	12'h0xd48: q<=8'b10010101;
	12'h0xd49: q<=8'b01100000;
	12'h0xd4a: q<=8'b10101001;
	12'h0xd4b: q<=8'b00000000;
	12'h0xd4c: q<=8'b11100101;
	12'h0xd4d: q<=8'b01011011;
	12'h0xd4e: q<=8'b10001101;
	12'h0xd4f: q<=8'b10010110;
	12'h0xd50: q<=8'b01100000;
	12'h0xd51: q<=8'b10101001;
	12'h0xd52: q<=8'b00011000;
	12'h0xd53: q<=8'b10001101;
	12'h0xd54: q<=8'b10001100;
	12'h0xd55: q<=8'b01100000;
	12'h0xd56: q<=8'b10100101;
	12'h0xd57: q<=8'b10100000;
	12'h0xd58: q<=8'b10001101;
	12'h0xd59: q<=8'b10001110;
	12'h0xd5a: q<=8'b01100000;
	12'h0xd5b: q<=8'b10001101;
	12'h0xd5c: q<=8'b10010100;
	12'h0xd5d: q<=8'b01100000;
	12'h0xd5e: q<=8'b00101100;
	12'h0xd5f: q<=8'b01000000;
	12'h0xd60: q<=8'b01100000;
	12'h0xd61: q<=8'b00110000;
	12'h0xd62: q<=8'b11111011;
	12'h0xd63: q<=8'b10101101;
	12'h0xd64: q<=8'b01100000;
	12'h0xd65: q<=8'b01100000;
	12'h0xd66: q<=8'b10000101;
	12'h0xd67: q<=8'b01111001;
	12'h0xd68: q<=8'b10101101;
	12'h0xd69: q<=8'b01110000;
	12'h0xd6a: q<=8'b01100000;
	12'h0xd6b: q<=8'b10000101;
	12'h0xd6c: q<=8'b01111010;
	12'h0xd6d: q<=8'b10100010;
	12'h0xd6e: q<=8'b00001111;
	12'h0xd6f: q<=8'b10001110;
	12'h0xd70: q<=8'b10001100;
	12'h0xd71: q<=8'b01100000;
	12'h0xd72: q<=8'b00111000;
	12'h0xd73: q<=8'b11101001;
	12'h0xd74: q<=8'b00000001;
	12'h0xd75: q<=8'b11010000;
	12'h0xd76: q<=8'b00000010;
	12'h0xd77: q<=8'b10101001;
	12'h0xd78: q<=8'b00000001;
	12'h0xd79: q<=8'b10100010;
	12'h0xd7a: q<=8'b00000000;
	12'h0xd7b: q<=8'b11101000;
	12'h0xd7c: q<=8'b00000110;
	12'h0xd7d: q<=8'b01111001;
	12'h0xd7e: q<=8'b00101010;
	12'h0xd7f: q<=8'b10010000;
	12'h0xd80: q<=8'b11111010;
	12'h0xd81: q<=8'b01001010;
	12'h0xd82: q<=8'b01001001;
	12'h0xd83: q<=8'b01111111;
	12'h0xd84: q<=8'b00011000;
	12'h0xd85: q<=8'b01101001;
	12'h0xd86: q<=8'b00000001;
	12'h0xd87: q<=8'b10101000;
	12'h0xd88: q<=8'b10001010;
	12'h0xd89: q<=8'b10111000;
	12'h0xd8a: q<=8'b01010000;
	12'h0xd8b: q<=8'b00000100;
	12'h0xd8c: q<=8'b10101001;
	12'h0xd8d: q<=8'b00000001;
	12'h0xd8e: q<=8'b10100000;
	12'h0xd8f: q<=8'b00000000;
	12'h0xd90: q<=8'b10000101;
	12'h0xd91: q<=8'b01111000;
	12'h0xd92: q<=8'b01001000;
	12'h0xd93: q<=8'b10011000;
	12'h0xd94: q<=8'b10100100;
	12'h0xd95: q<=8'b10101001;
	12'h0xd96: q<=8'b10010001;
	12'h0xd97: q<=8'b01110100;
	12'h0xd98: q<=8'b11001000;
	12'h0xd99: q<=8'b01101000;
	12'h0xd9a: q<=8'b00001001;
	12'h0xd9b: q<=8'b01110000;
	12'h0xd9c: q<=8'b10010001;
	12'h0xd9d: q<=8'b01110100;
	12'h0xd9e: q<=8'b11001000;
	12'h0xd9f: q<=8'b01100000;
	12'h0xda0: q<=8'b10000101;
	12'h0xda1: q<=8'b00110110;
	12'h0xda2: q<=8'b10111001;
	12'h0xda3: q<=8'b11001110;
	12'h0xda4: q<=8'b00000011;
	12'h0xda5: q<=8'b10000101;
	12'h0xda6: q<=8'b01010110;
	12'h0xda7: q<=8'b10111001;
	12'h0xda8: q<=8'b11011110;
	12'h0xda9: q<=8'b00000011;
	12'h0xdaa: q<=8'b10000101;
	12'h0xdab: q<=8'b01011000;
	12'h0xdac: q<=8'b10100101;
	12'h0xdad: q<=8'b01010111;
	12'h0xdae: q<=8'b10000101;
	12'h0xdaf: q<=8'b00101111;
	12'h0xdb0: q<=8'b10011000;
	12'h0xdb1: q<=8'b00011000;
	12'h0xdb2: q<=8'b01101001;
	12'h0xdb3: q<=8'b00000001;
	12'h0xdb4: q<=8'b00101001;
	12'h0xdb5: q<=8'b00001111;
	12'h0xdb6: q<=8'b10101010;
	12'h0xdb7: q<=8'b10111101;
	12'h0xdb8: q<=8'b11001110;
	12'h0xdb9: q<=8'b00000011;
	12'h0xdba: q<=8'b10000101;
	12'h0xdbb: q<=8'b00101110;
	12'h0xdbc: q<=8'b10111101;
	12'h0xdbd: q<=8'b11011110;
	12'h0xdbe: q<=8'b00000011;
	12'h0xdbf: q<=8'b10000101;
	12'h0xdc0: q<=8'b00110000;
	12'h0xdc1: q<=8'b10101001;
	12'h0xdc2: q<=8'b00000000;
	12'h0xdc3: q<=8'b10000101;
	12'h0xdc4: q<=8'b01011001;
	12'h0xdc5: q<=8'b10101001;
	12'h0xdc6: q<=8'b00000100;
	12'h0xdc7: q<=8'b10000101;
	12'h0xdc8: q<=8'b01011010;
	12'h0xdc9: q<=8'b10100100;
	12'h0xdca: q<=8'b00110110;
	12'h0xdcb: q<=8'b10100101;
	12'h0xdcc: q<=8'b01011011;
	12'h0xdcd: q<=8'b00110000;
	12'h0xdce: q<=8'b00000111;
	12'h0xdcf: q<=8'b10100101;
	12'h0xdd0: q<=8'b01010111;
	12'h0xdd1: q<=8'b11000101;
	12'h0xdd2: q<=8'b01011111;
	12'h0xdd3: q<=8'b10110000;
	12'h0xdd4: q<=8'b00000001;
	12'h0xdd5: q<=8'b01100000;
	12'h0xdd6: q<=8'b10111001;
	12'h0xdd7: q<=8'b10110110;
	12'h0xdd8: q<=8'b10111111;
	12'h0xdd9: q<=8'b10000101;
	12'h0xdda: q<=8'b10011001;
	12'h0xddb: q<=8'b10111001;
	12'h0xddc: q<=8'b11000100;
	12'h0xddd: q<=8'b10111111;
	12'h0xdde: q<=8'b10000101;
	12'h0xddf: q<=8'b00111000;
	12'h0xde0: q<=8'b10100100;
	12'h0xde1: q<=8'b10011110;
	12'h0xde2: q<=8'b10101001;
	12'h0xde3: q<=8'b00001000;
	12'h0xde4: q<=8'b00100000;
	12'h0xde5: q<=8'b01001100;
	12'h0xde6: q<=8'b11011111;
	12'h0xde7: q<=8'b00100000;
	12'h0xde8: q<=8'b10011000;
	12'h0xde9: q<=8'b11000000;
	12'h0xdea: q<=8'b10100010;
	12'h0xdeb: q<=8'b01100001;
	12'h0xdec: q<=8'b00100000;
	12'h0xded: q<=8'b01100101;
	12'h0xdee: q<=8'b11000111;
	12'h0xdef: q<=8'b10100101;
	12'h0xdf0: q<=8'b00101110;
	12'h0xdf1: q<=8'b10000101;
	12'h0xdf2: q<=8'b01010110;
	12'h0xdf3: q<=8'b10100101;
	12'h0xdf4: q<=8'b00101111;
	12'h0xdf5: q<=8'b10000101;
	12'h0xdf6: q<=8'b01010111;
	12'h0xdf7: q<=8'b10100101;
	12'h0xdf8: q<=8'b00110000;
	12'h0xdf9: q<=8'b10000101;
	12'h0xdfa: q<=8'b01011000;
	12'h0xdfb: q<=8'b00100000;
	12'h0xdfc: q<=8'b10011000;
	12'h0xdfd: q<=8'b11000000;
	12'h0xdfe: q<=8'b10100100;
	12'h0xdff: q<=8'b01011001;
	12'h0xe00: q<=8'b10100101;
	12'h0xe01: q<=8'b01011010;
	12'h0xe02: q<=8'b00100000;
	12'h0xe03: q<=8'b01101100;
	12'h0xe04: q<=8'b11011111;
	12'h0xe05: q<=8'b10100101;
	12'h0xe06: q<=8'b01100001;
	12'h0xe07: q<=8'b00111000;
	12'h0xe08: q<=8'b11100101;
	12'h0xe09: q<=8'b01101010;
	12'h0xe0a: q<=8'b10000101;
	12'h0xe0b: q<=8'b01111001;
	12'h0xe0c: q<=8'b10100101;
	12'h0xe0d: q<=8'b01100010;
	12'h0xe0e: q<=8'b11100101;
	12'h0xe0f: q<=8'b01101011;
	12'h0xe10: q<=8'b10000101;
	12'h0xe11: q<=8'b10011011;
	12'h0xe12: q<=8'b00110000;
	12'h0xe13: q<=8'b00001001;
	12'h0xe14: q<=8'b11110000;
	12'h0xe15: q<=8'b00000100;
	12'h0xe16: q<=8'b10101001;
	12'h0xe17: q<=8'b11111111;
	12'h0xe18: q<=8'b10000101;
	12'h0xe19: q<=8'b01111001;
	12'h0xe1a: q<=8'b10111000;
	12'h0xe1b: q<=8'b01010000;
	12'h0xe1c: q<=8'b00010110;
	12'h0xe1d: q<=8'b11001001;
	12'h0xe1e: q<=8'b11111111;
	12'h0xe1f: q<=8'b11110000;
	12'h0xe20: q<=8'b00000101;
	12'h0xe21: q<=8'b10101001;
	12'h0xe22: q<=8'b11111111;
	12'h0xe23: q<=8'b10111000;
	12'h0xe24: q<=8'b01010000;
	12'h0xe25: q<=8'b00001011;
	12'h0xe26: q<=8'b10100101;
	12'h0xe27: q<=8'b01111001;
	12'h0xe28: q<=8'b01001001;
	12'h0xe29: q<=8'b11111111;
	12'h0xe2a: q<=8'b00011000;
	12'h0xe2b: q<=8'b01101001;
	12'h0xe2c: q<=8'b00000001;
	12'h0xe2d: q<=8'b10010000;
	12'h0xe2e: q<=8'b00000010;
	12'h0xe2f: q<=8'b10101001;
	12'h0xe30: q<=8'b11111111;
	12'h0xe31: q<=8'b10000101;
	12'h0xe32: q<=8'b01111001;
	12'h0xe33: q<=8'b10100101;
	12'h0xe34: q<=8'b01100011;
	12'h0xe35: q<=8'b00111000;
	12'h0xe36: q<=8'b11100101;
	12'h0xe37: q<=8'b01101100;
	12'h0xe38: q<=8'b10000101;
	12'h0xe39: q<=8'b10001001;
	12'h0xe3a: q<=8'b10100101;
	12'h0xe3b: q<=8'b01100100;
	12'h0xe3c: q<=8'b11100101;
	12'h0xe3d: q<=8'b01101101;
	12'h0xe3e: q<=8'b10000101;
	12'h0xe3f: q<=8'b10011101;
	12'h0xe40: q<=8'b00110000;
	12'h0xe41: q<=8'b00001001;
	12'h0xe42: q<=8'b11110000;
	12'h0xe43: q<=8'b00000100;
	12'h0xe44: q<=8'b10101001;
	12'h0xe45: q<=8'b11111111;
	12'h0xe46: q<=8'b10000101;
	12'h0xe47: q<=8'b10001001;
	12'h0xe48: q<=8'b10111000;
	12'h0xe49: q<=8'b01010000;
	12'h0xe4a: q<=8'b00010010;
	12'h0xe4b: q<=8'b11001001;
	12'h0xe4c: q<=8'b11111111;
	12'h0xe4d: q<=8'b11110000;
	12'h0xe4e: q<=8'b00000101;
	12'h0xe4f: q<=8'b10101001;
	12'h0xe50: q<=8'b11111111;
	12'h0xe51: q<=8'b10111000;
	12'h0xe52: q<=8'b01010000;
	12'h0xe53: q<=8'b00000111;
	12'h0xe54: q<=8'b10100101;
	12'h0xe55: q<=8'b10001001;
	12'h0xe56: q<=8'b01001001;
	12'h0xe57: q<=8'b11111111;
	12'h0xe58: q<=8'b00011000;
	12'h0xe59: q<=8'b01101001;
	12'h0xe5a: q<=8'b00000001;
	12'h0xe5b: q<=8'b10000101;
	12'h0xe5c: q<=8'b10001001;
	12'h0xe5d: q<=8'b10101001;
	12'h0xe5e: q<=8'b00000000;
	12'h0xe5f: q<=8'b10000101;
	12'h0xe60: q<=8'b10000010;
	12'h0xe61: q<=8'b10000101;
	12'h0xe62: q<=8'b10010010;
	12'h0xe63: q<=8'b10100101;
	12'h0xe64: q<=8'b01111001;
	12'h0xe65: q<=8'b00001010;
	12'h0xe66: q<=8'b00100110;
	12'h0xe67: q<=8'b10000010;
	12'h0xe68: q<=8'b10000101;
	12'h0xe69: q<=8'b01111010;
	12'h0xe6a: q<=8'b00001010;
	12'h0xe6b: q<=8'b10000101;
	12'h0xe6c: q<=8'b01111100;
	12'h0xe6d: q<=8'b10100101;
	12'h0xe6e: q<=8'b10000010;
	12'h0xe6f: q<=8'b00101010;
	12'h0xe70: q<=8'b10000101;
	12'h0xe71: q<=8'b10000100;
	12'h0xe72: q<=8'b10100101;
	12'h0xe73: q<=8'b01111100;
	12'h0xe74: q<=8'b01100101;
	12'h0xe75: q<=8'b01111001;
	12'h0xe76: q<=8'b10000101;
	12'h0xe77: q<=8'b01111101;
	12'h0xe78: q<=8'b10100101;
	12'h0xe79: q<=8'b10000100;
	12'h0xe7a: q<=8'b01101001;
	12'h0xe7b: q<=8'b00000000;
	12'h0xe7c: q<=8'b10000101;
	12'h0xe7d: q<=8'b10000101;
	12'h0xe7e: q<=8'b10100101;
	12'h0xe7f: q<=8'b01111010;
	12'h0xe80: q<=8'b01100101;
	12'h0xe81: q<=8'b01111001;
	12'h0xe82: q<=8'b10000101;
	12'h0xe83: q<=8'b01111011;
	12'h0xe84: q<=8'b10100101;
	12'h0xe85: q<=8'b10000010;
	12'h0xe86: q<=8'b01101001;
	12'h0xe87: q<=8'b00000000;
	12'h0xe88: q<=8'b10000101;
	12'h0xe89: q<=8'b10000011;
	12'h0xe8a: q<=8'b10000101;
	12'h0xe8b: q<=8'b10000110;
	12'h0xe8c: q<=8'b10100101;
	12'h0xe8d: q<=8'b01111011;
	12'h0xe8e: q<=8'b00001010;
	12'h0xe8f: q<=8'b10000101;
	12'h0xe90: q<=8'b01111110;
	12'h0xe91: q<=8'b00100110;
	12'h0xe92: q<=8'b10000110;
	12'h0xe93: q<=8'b01100101;
	12'h0xe94: q<=8'b01111001;
	12'h0xe95: q<=8'b10000101;
	12'h0xe96: q<=8'b01111111;
	12'h0xe97: q<=8'b10100101;
	12'h0xe98: q<=8'b10000110;
	12'h0xe99: q<=8'b01101001;
	12'h0xe9a: q<=8'b00000000;
	12'h0xe9b: q<=8'b10000101;
	12'h0xe9c: q<=8'b10000111;
	12'h0xe9d: q<=8'b10100101;
	12'h0xe9e: q<=8'b10001001;
	12'h0xe9f: q<=8'b00001010;
	12'h0xea0: q<=8'b00100110;
	12'h0xea1: q<=8'b10010010;
	12'h0xea2: q<=8'b10000101;
	12'h0xea3: q<=8'b10001010;
	12'h0xea4: q<=8'b00001010;
	12'h0xea5: q<=8'b10000101;
	12'h0xea6: q<=8'b10001100;
	12'h0xea7: q<=8'b10100101;
	12'h0xea8: q<=8'b10010010;
	12'h0xea9: q<=8'b00101010;
	12'h0xeaa: q<=8'b10000101;
	12'h0xeab: q<=8'b10010100;
	12'h0xeac: q<=8'b10100101;
	12'h0xead: q<=8'b10001100;
	12'h0xeae: q<=8'b01100101;
	12'h0xeaf: q<=8'b10001001;
	12'h0xeb0: q<=8'b10000101;
	12'h0xeb1: q<=8'b10001101;
	12'h0xeb2: q<=8'b10100101;
	12'h0xeb3: q<=8'b10010100;
	12'h0xeb4: q<=8'b01101001;
	12'h0xeb5: q<=8'b00000000;
	12'h0xeb6: q<=8'b10000101;
	12'h0xeb7: q<=8'b10010101;
	12'h0xeb8: q<=8'b10100101;
	12'h0xeb9: q<=8'b10001010;
	12'h0xeba: q<=8'b01100101;
	12'h0xebb: q<=8'b10001001;
	12'h0xebc: q<=8'b10000101;
	12'h0xebd: q<=8'b10001011;
	12'h0xebe: q<=8'b10100101;
	12'h0xebf: q<=8'b10010010;
	12'h0xec0: q<=8'b01101001;
	12'h0xec1: q<=8'b00000000;
	12'h0xec2: q<=8'b10000101;
	12'h0xec3: q<=8'b10010011;
	12'h0xec4: q<=8'b10000101;
	12'h0xec5: q<=8'b10010110;
	12'h0xec6: q<=8'b10100101;
	12'h0xec7: q<=8'b10001011;
	12'h0xec8: q<=8'b00001010;
	12'h0xec9: q<=8'b10000101;
	12'h0xeca: q<=8'b10001110;
	12'h0xecb: q<=8'b00100110;
	12'h0xecc: q<=8'b10010110;
	12'h0xecd: q<=8'b01100101;
	12'h0xece: q<=8'b10001001;
	12'h0xecf: q<=8'b10000101;
	12'h0xed0: q<=8'b10001111;
	12'h0xed1: q<=8'b10100101;
	12'h0xed2: q<=8'b10010110;
	12'h0xed3: q<=8'b01101001;
	12'h0xed4: q<=8'b00000000;
	12'h0xed5: q<=8'b10000101;
	12'h0xed6: q<=8'b10010111;
	12'h0xed7: q<=8'b10100000;
	12'h0xed8: q<=8'b00000000;
	12'h0xed9: q<=8'b10000100;
	12'h0xeda: q<=8'b10101001;
	12'h0xedb: q<=8'b10100100;
	12'h0xedc: q<=8'b00111000;
	12'h0xedd: q<=8'b10111001;
	12'h0xede: q<=8'b11010011;
	12'h0xedf: q<=8'b10111111;
	12'h0xee0: q<=8'b11001001;
	12'h0xee1: q<=8'b00000001;
	12'h0xee2: q<=8'b11010000;
	12'h0xee3: q<=8'b00000010;
	12'h0xee4: q<=8'b10101001;
	12'h0xee5: q<=8'b11000000;
	12'h0xee6: q<=8'b10000101;
	12'h0xee7: q<=8'b01110011;
	12'h0xee8: q<=8'b10111001;
	12'h0xee9: q<=8'b11010010;
	12'h0xeea: q<=8'b10111111;
	12'h0xeeb: q<=8'b10000101;
	12'h0xeec: q<=8'b00101101;
	12'h0xeed: q<=8'b11001000;
	12'h0xeee: q<=8'b11001000;
	12'h0xeef: q<=8'b10000100;
	12'h0xef0: q<=8'b00111000;
	12'h0xef1: q<=8'b10101010;
	12'h0xef2: q<=8'b00101001;
	12'h0xef3: q<=8'b00000111;
	12'h0xef4: q<=8'b10101000;
	12'h0xef5: q<=8'b10001010;
	12'h0xef6: q<=8'b00001010;
	12'h0xef7: q<=8'b10000101;
	12'h0xef8: q<=8'b00101011;
	12'h0xef9: q<=8'b01001010;
	12'h0xefa: q<=8'b01001010;
	12'h0xefb: q<=8'b01001010;
	12'h0xefc: q<=8'b01001010;
	12'h0xefd: q<=8'b00101001;
	12'h0xefe: q<=8'b00000111;
	12'h0xeff: q<=8'b10101010;
	12'h0xf00: q<=8'b10100101;
	12'h0xf01: q<=8'b00101011;
	12'h0xf02: q<=8'b01000101;
	12'h0xf03: q<=8'b10011011;
	12'h0xf04: q<=8'b00110000;
	12'h0xf05: q<=8'b00001011;
	12'h0xf06: q<=8'b10111001;
	12'h0xf07: q<=8'b01111000;
	12'h0xf08: q<=8'b00000000;
	12'h0xf09: q<=8'b10000101;
	12'h0xf0a: q<=8'b01100001;
	12'h0xf0b: q<=8'b10111001;
	12'h0xf0c: q<=8'b10000000;
	12'h0xf0d: q<=8'b00000000;
	12'h0xf0e: q<=8'b10111000;
	12'h0xf0f: q<=8'b01010000;
	12'h0xf10: q<=8'b00010001;
	12'h0xf11: q<=8'b10111001;
	12'h0xf12: q<=8'b01111000;
	12'h0xf13: q<=8'b00000000;
	12'h0xf14: q<=8'b01001001;
	12'h0xf15: q<=8'b11111111;
	12'h0xf16: q<=8'b00011000;
	12'h0xf17: q<=8'b01101001;
	12'h0xf18: q<=8'b00000001;
	12'h0xf19: q<=8'b10000101;
	12'h0xf1a: q<=8'b01100001;
	12'h0xf1b: q<=8'b10111001;
	12'h0xf1c: q<=8'b10000000;
	12'h0xf1d: q<=8'b00000000;
	12'h0xf1e: q<=8'b01001001;
	12'h0xf1f: q<=8'b11111111;
	12'h0xf20: q<=8'b01101001;
	12'h0xf21: q<=8'b00000000;
	12'h0xf22: q<=8'b10000101;
	12'h0xf23: q<=8'b01100010;
	12'h0xf24: q<=8'b10100101;
	12'h0xf25: q<=8'b00101101;
	12'h0xf26: q<=8'b01000101;
	12'h0xf27: q<=8'b10011101;
	12'h0xf28: q<=8'b00010000;
	12'h0xf29: q<=8'b00001110;
	12'h0xf2a: q<=8'b10110101;
	12'h0xf2b: q<=8'b10001000;
	12'h0xf2c: q<=8'b00011000;
	12'h0xf2d: q<=8'b01100101;
	12'h0xf2e: q<=8'b01100001;
	12'h0xf2f: q<=8'b10000101;
	12'h0xf30: q<=8'b01100001;
	12'h0xf31: q<=8'b10110101;
	12'h0xf32: q<=8'b10010000;
	12'h0xf33: q<=8'b01100101;
	12'h0xf34: q<=8'b01100010;
	12'h0xf35: q<=8'b10111000;
	12'h0xf36: q<=8'b01010000;
	12'h0xf37: q<=8'b00001011;
	12'h0xf38: q<=8'b10100101;
	12'h0xf39: q<=8'b01100001;
	12'h0xf3a: q<=8'b00111000;
	12'h0xf3b: q<=8'b11110101;
	12'h0xf3c: q<=8'b10001000;
	12'h0xf3d: q<=8'b10000101;
	12'h0xf3e: q<=8'b01100001;
	12'h0xf3f: q<=8'b10100101;
	12'h0xf40: q<=8'b01100010;
	12'h0xf41: q<=8'b11110101;
	12'h0xf42: q<=8'b10010000;
	12'h0xf43: q<=8'b10000101;
	12'h0xf44: q<=8'b01100010;
	12'h0xf45: q<=8'b10100101;
	12'h0xf46: q<=8'b00101011;
	12'h0xf47: q<=8'b01000101;
	12'h0xf48: q<=8'b10011101;
	12'h0xf49: q<=8'b00110000;
	12'h0xf4a: q<=8'b00001011;
	12'h0xf4b: q<=8'b10111001;
	12'h0xf4c: q<=8'b10001000;
	12'h0xf4d: q<=8'b00000000;
	12'h0xf4e: q<=8'b10000101;
	12'h0xf4f: q<=8'b01100011;
	12'h0xf50: q<=8'b10111001;
	12'h0xf51: q<=8'b10010000;
	12'h0xf52: q<=8'b00000000;
	12'h0xf53: q<=8'b10111000;
	12'h0xf54: q<=8'b01010000;
	12'h0xf55: q<=8'b00010001;
	12'h0xf56: q<=8'b10111001;
	12'h0xf57: q<=8'b10001000;
	12'h0xf58: q<=8'b00000000;
	12'h0xf59: q<=8'b01001001;
	12'h0xf5a: q<=8'b11111111;
	12'h0xf5b: q<=8'b00011000;
	12'h0xf5c: q<=8'b01101001;
	12'h0xf5d: q<=8'b00000001;
	12'h0xf5e: q<=8'b10000101;
	12'h0xf5f: q<=8'b01100011;
	12'h0xf60: q<=8'b10111001;
	12'h0xf61: q<=8'b10010000;
	12'h0xf62: q<=8'b00000000;
	12'h0xf63: q<=8'b01001001;
	12'h0xf64: q<=8'b11111111;
	12'h0xf65: q<=8'b01101001;
	12'h0xf66: q<=8'b00000000;
	12'h0xf67: q<=8'b10000101;
	12'h0xf68: q<=8'b01100100;
	12'h0xf69: q<=8'b10100101;
	12'h0xf6a: q<=8'b00101101;
	12'h0xf6b: q<=8'b01000101;
	12'h0xf6c: q<=8'b10011011;
	12'h0xf6d: q<=8'b00010000;
	12'h0xf6e: q<=8'b00001110;
	12'h0xf6f: q<=8'b10100101;
	12'h0xf70: q<=8'b01100011;
	12'h0xf71: q<=8'b00111000;
	12'h0xf72: q<=8'b11110101;
	12'h0xf73: q<=8'b01111000;
	12'h0xf74: q<=8'b10000101;
	12'h0xf75: q<=8'b01100011;
	12'h0xf76: q<=8'b10100101;
	12'h0xf77: q<=8'b01100100;
	12'h0xf78: q<=8'b11110101;
	12'h0xf79: q<=8'b10000000;
	12'h0xf7a: q<=8'b10111000;
	12'h0xf7b: q<=8'b01010000;
	12'h0xf7c: q<=8'b00001011;
	12'h0xf7d: q<=8'b10100101;
	12'h0xf7e: q<=8'b01100011;
	12'h0xf7f: q<=8'b00011000;
	12'h0xf80: q<=8'b01110101;
	12'h0xf81: q<=8'b01111000;
	12'h0xf82: q<=8'b10000101;
	12'h0xf83: q<=8'b01100011;
	12'h0xf84: q<=8'b10100101;
	12'h0xf85: q<=8'b01100100;
	12'h0xf86: q<=8'b01110101;
	12'h0xf87: q<=8'b10000000;
	12'h0xf88: q<=8'b10000101;
	12'h0xf89: q<=8'b01100100;
	12'h0xf8a: q<=8'b10100100;
	12'h0xf8b: q<=8'b10101001;
	12'h0xf8c: q<=8'b10100101;
	12'h0xf8d: q<=8'b01100011;
	12'h0xf8e: q<=8'b10010001;
	12'h0xf8f: q<=8'b01110100;
	12'h0xf90: q<=8'b11001000;
	12'h0xf91: q<=8'b10100101;
	12'h0xf92: q<=8'b01100100;
	12'h0xf93: q<=8'b00101001;
	12'h0xf94: q<=8'b00011111;
	12'h0xf95: q<=8'b10010001;
	12'h0xf96: q<=8'b01110100;
	12'h0xf97: q<=8'b11001000;
	12'h0xf98: q<=8'b10100101;
	12'h0xf99: q<=8'b01100001;
	12'h0xf9a: q<=8'b10010001;
	12'h0xf9b: q<=8'b01110100;
	12'h0xf9c: q<=8'b11001000;
	12'h0xf9d: q<=8'b10100101;
	12'h0xf9e: q<=8'b01100010;
	12'h0xf9f: q<=8'b00101001;
	12'h0xfa0: q<=8'b00011111;
	12'h0xfa1: q<=8'b00000101;
	12'h0xfa2: q<=8'b01110011;
	12'h0xfa3: q<=8'b10010001;
	12'h0xfa4: q<=8'b01110100;
	12'h0xfa5: q<=8'b11001000;
	12'h0xfa6: q<=8'b10000100;
	12'h0xfa7: q<=8'b10101001;
	12'h0xfa8: q<=8'b11000110;
	12'h0xfa9: q<=8'b10011001;
	12'h0xfaa: q<=8'b11110000;
	12'h0xfab: q<=8'b00000011;
	12'h0xfac: q<=8'b01001100;
	12'h0xfad: q<=8'b11011011;
	12'h0xfae: q<=8'b10111110;
	12'h0xfaf: q<=8'b10100100;
	12'h0xfb0: q<=8'b10101001;
	12'h0xfb1: q<=8'b10001000;
	12'h0xfb2: q<=8'b01001100;
	12'h0xfb3: q<=8'b01011111;
	12'h0xfb4: q<=8'b11011111;
	12'h0xfb5: q<=8'b00001000;
	12'h0xfb6: q<=8'b00001000;
	12'h0xfb7: q<=8'b00001000;
	12'h0xfb8: q<=8'b00001000;
	12'h0xfb9: q<=8'b00001000;
	12'h0xfba: q<=8'b00001000;
	12'h0xfbb: q<=8'b00001000;
	12'h0xfbc: q<=8'b00001000;
	12'h0xfbd: q<=8'b00001000;
	12'h0xfbe: q<=8'b00001001;
	12'h0xfbf: q<=8'b00000110;
	12'h0xfc0: q<=8'b00000111;
	12'h0xfc1: q<=8'b00000111;
	12'h0xfc2: q<=8'b00000100;
	12'h0xfc3: q<=8'b00000010;
	12'h0xfc4: q<=8'b00000000;
	12'h0xfc5: q<=8'b00010000;
	12'h0xfc6: q<=8'b00100000;
	12'h0xfc7: q<=8'b00110000;
	12'h0xfc8: q<=8'b01000000;
	12'h0xfc9: q<=8'b01010000;
	12'h0xfca: q<=8'b01100000;
	12'h0xfcb: q<=8'b01110000;
	12'h0xfcc: q<=8'b10000000;
	12'h0xfcd: q<=8'b10010010;
	12'h0xfce: q<=8'b10011110;
	12'h0xfcf: q<=8'b10101100;
	12'h0xfd0: q<=8'b10111010;
	12'h0xfd1: q<=8'b11000010;
	12'h0xfd2: q<=8'b00001100;
	12'h0xfd3: q<=8'b00000001;
	12'h0xfd4: q<=8'b10001100;
	12'h0xfd5: q<=8'b00000001;
	12'h0xfd6: q<=8'b01001010;
	12'h0xfd7: q<=8'b00000001;
	12'h0xfd8: q<=8'b00001001;
	12'h0xfd9: q<=8'b00000001;
	12'h0xfda: q<=8'b11001011;
	12'h0xfdb: q<=8'b00000001;
	12'h0xfdc: q<=8'b01001011;
	12'h0xfdd: q<=8'b00000001;
	12'h0xfde: q<=8'b10001001;
	12'h0xfdf: q<=8'b00000001;
	12'h0xfe0: q<=8'b11001010;
	12'h0xfe1: q<=8'b00000001;
	12'h0xfe2: q<=8'b10010000;
	12'h0xfe3: q<=8'b00000001;
	12'h0xfe4: q<=8'b10001010;
	12'h0xfe5: q<=8'b00000001;
	12'h0xfe6: q<=8'b00100011;
	12'h0xfe7: q<=8'b00000001;
	12'h0xfe8: q<=8'b11011011;
	12'h0xfe9: q<=8'b00000001;
	12'h0xfea: q<=8'b01000001;
	12'h0xfeb: q<=8'b00000001;
	12'h0xfec: q<=8'b00010000;
	12'h0xfed: q<=8'b00000001;
	12'h0xfee: q<=8'b00001010;
	12'h0xfef: q<=8'b00000001;
	12'h0xff0: q<=8'b11001011;
	12'h0xff1: q<=8'b00000001;
	12'h0xff2: q<=8'b10010001;
	12'h0xff3: q<=8'b00000001;
	12'h0xff4: q<=8'b00010111;
	12'h0xff5: q<=8'b00000001;
	12'h0xff6: q<=8'b01001011;
	12'h0xff7: q<=8'b00000001;
	12'h0xff8: q<=8'b10001010;
	12'h0xff9: q<=8'b00000001;
	12'h0xffa: q<=8'b11001110;
	12'h0xffb: q<=8'b00000001;
	12'h0xffc: q<=8'b00001000;
	12'h0xffd: q<=8'b00000001;
	12'h0xffe: q<=8'b00001010;
	12'h0xfff: q<=8'b00000001;
endcase
end
assign dout=q;
endmodule
