module rom_CombinedROM
(
input clk,
input [7:0] addr,
output [23:0] dout,
input cs );
reg [23:0] q;
always @(posedge clk) 
begin 
case (addr) 
	8'h0x0: q<=24'b000000000001011100000000;
	8'h0x1: q<=24'b000000010010000010011100;
	8'h0x2: q<=24'b000001000010001010011101;
	8'h0x3: q<=24'b000000110010100010010100;
	8'h0x4: q<=24'b000000000010000000110000;
	8'h0x5: q<=24'b000000010100010000110000;
	8'h0x6: q<=24'b000000000010010000000000;
	8'h0x7: q<=24'b000100010001000001001000;
	8'h0x8: q<=24'b000000010001000001000010;
	8'h0x9: q<=24'b000001110010000010011100;
	8'h0xa: q<=24'b000000010011000001100000;
	8'h0xb: q<=24'b000011010010001010011101;
	8'h0xc: q<=24'b000011000010100010010100;
	8'h0xd: q<=24'b000010100000000010010000;
	8'h0xe: q<=24'b000000010011000000011100;
	8'h0xf: q<=24'b000001110000000010010100;
	8'h0x10: q<=24'b000000000011101100010000;
	8'h0x11: q<=24'b000000010011101100010000;
	8'h0x12: q<=24'b000000100011101100010000;
	8'h0x13: q<=24'b000000110011101100010000;
	8'h0x14: q<=24'b000001000011101100010000;
	8'h0x15: q<=24'b000001010011101100010000;
	8'h0x16: q<=24'b101110110010010010000100;
	8'h0x17: q<=24'b000001110011101100010000;
	8'h0x18: q<=24'b000010000011101100010000;
	8'h0x19: q<=24'b000010010011101100010000;
	8'h0x1a: q<=24'b000010100011101100010000;
	8'h0x1b: q<=24'b000010110011101100010000;
	8'h0x1c: q<=24'b000011000011101100010000;
	8'h0x1d: q<=24'b000011010011101100010000;
	8'h0x1e: q<=24'b000011100011101100010000;
	8'h0x1f: q<=24'b000011110011101100010000;
	8'h0x20: q<=24'b000100000111001110110100;
	8'h0x21: q<=24'b000100001011001110110100;
	8'h0x22: q<=24'b000100010111001110110100;
	8'h0x23: q<=24'b000100011011001110110100;
	8'h0x24: q<=24'b000100100111001110110100;
	8'h0x25: q<=24'b000100101011001110110100;
	8'h0x26: q<=24'b000100110111001110110100;
	8'h0x27: q<=24'b000100111011001110110100;
	8'h0x28: q<=24'b000101000111001110110100;
	8'h0x29: q<=24'b000101001011001110110100;
	8'h0x2a: q<=24'b000101010111001110110100;
	8'h0x2b: q<=24'b000101011011001110110100;
	8'h0x2c: q<=24'b000101100111001110110100;
	8'h0x2d: q<=24'b000101101011001110110100;
	8'h0x2e: q<=24'b000101110111001110110100;
	8'h0x2f: q<=24'b000101111011001110110100;
	8'h0x30: q<=24'b000110000111001110110100;
	8'h0x31: q<=24'b000110001011001110110100;
	8'h0x32: q<=24'b000110010111001110110100;
	8'h0x33: q<=24'b000110011011001110110100;
	8'h0x34: q<=24'b000110100111001110110100;
	8'h0x35: q<=24'b000110101011001110110100;
	8'h0x36: q<=24'b000110110111001110110100;
	8'h0x37: q<=24'b000110111011001110110100;
	8'h0x38: q<=24'b000111000111001110110100;
	8'h0x39: q<=24'b000111001011001110110100;
	8'h0x3a: q<=24'b000111010111001110110100;
	8'h0x3b: q<=24'b000111011011001110110100;
	8'h0x3c: q<=24'b000111100111001110110100;
	8'h0x3d: q<=24'b000111101011001110110100;
	8'h0x3e: q<=24'b000111110111001110110100;
	8'h0x3f: q<=24'b000111111011001110110100;
	8'h0x40: q<=24'b000000000010101100010000;
	8'h0x41: q<=24'b010001011011001110110100;
	8'h0x42: q<=24'b000001011011001100110000;
	8'h0x43: q<=24'b000011110011010000110000;
	8'h0x44: q<=24'b010010000000000010010100;
	8'h0x45: q<=24'b111111110001011100110000;
	8'h0x46: q<=24'b001001000001000100110001;
	8'h0x47: q<=24'b001101010001000100110001;
	8'h0x48: q<=24'b000011011100000000110000;
	8'h0x49: q<=24'b010011001100000010001100;
	8'h0x4a: q<=24'b000000000010001000000001;
	8'h0x4b: q<=24'b000011010011001000110001;
	8'h0x4c: q<=24'b110011000001000101000001;
	8'h0x4d: q<=24'b110111000001000001001010;
	8'h0x4e: q<=24'b110111000001000001001010;
	8'h0x4f: q<=24'b110111000001000001001010;
	8'h0x50: q<=24'b110111000001000001001010;
	8'h0x51: q<=24'b110111000001000001001010;
	8'h0x52: q<=24'b110111000001000001001010;
	8'h0x53: q<=24'b110111000001000001001010;
	8'h0x54: q<=24'b110111000001000001001010;
	8'h0x55: q<=24'b110111000001000001001010;
	8'h0x56: q<=24'b110111000001000001001010;
	8'h0x57: q<=24'b110111000001000001001010;
	8'h0x58: q<=24'b110111000001000001001010;
	8'h0x59: q<=24'b110111000001000001001010;
	8'h0x5a: q<=24'b110111000001000001001010;
	8'h0x5b: q<=24'b110111000001000001001010;
	8'h0x5c: q<=24'b110111000001000001001010;
	8'h0x5d: q<=24'b000011100010000000110000;
	8'h0x5e: q<=24'b000111011100001000110001;
	8'h0x5f: q<=24'b011000110000000010010000;
	8'h0x60: q<=24'b000001010011000000001100;
	8'h0x61: q<=24'b000000000010001000000001;
	8'h0x62: q<=24'b000011010011001000110001;
	8'h0x63: q<=24'b011101110001000101000001;
	8'h0x64: q<=24'b110101110001000001001010;
	8'h0x65: q<=24'b110101110001000001001010;
	8'h0x66: q<=24'b110101110001000001001010;
	8'h0x67: q<=24'b110101110001000001001010;
	8'h0x68: q<=24'b110101110001000001001010;
	8'h0x69: q<=24'b110101110001000001001010;
	8'h0x6a: q<=24'b110101110001000001001010;
	8'h0x6b: q<=24'b110101110001000001001010;
	8'h0x6c: q<=24'b110101110001000001001010;
	8'h0x6d: q<=24'b110101110001000001001010;
	8'h0x6e: q<=24'b110101110001000001001010;
	8'h0x6f: q<=24'b110101110001000001001010;
	8'h0x70: q<=24'b110101110001000001001010;
	8'h0x71: q<=24'b110101110001000001001010;
	8'h0x72: q<=24'b110101110001000001001010;
	8'h0x73: q<=24'b110101110001000001001010;
	8'h0x74: q<=24'b110001110001000000110000;
	8'h0x75: q<=24'b000011100011000001010000;
	8'h0x76: q<=24'b000011000010000001010000;
	8'h0x77: q<=24'b110011100001000000000000;
	8'h0x78: q<=24'b011110100010000010011100;
	8'h0x79: q<=24'b000001110011000000110001;
	8'h0x7a: q<=24'b011111010000000010010000;
	8'h0x7b: q<=24'b000011110011000000011100;
	8'h0x7c: q<=24'b000001110011100000010000;
	8'h0x7d: q<=24'b001001110001000000110000;
	8'h0x7e: q<=24'b000111011100000000110000;
	8'h0x7f: q<=24'b100000110000000010010000;
	8'h0x80: q<=24'b000001000011000000001100;
	8'h0x81: q<=24'b000000000010001000000001;
	8'h0x82: q<=24'b110111010011001000110001;
	8'h0x83: q<=24'b110011000001000101000001;
	8'h0x84: q<=24'b110111000001000001001010;
	8'h0x85: q<=24'b110111000001000001001010;
	8'h0x86: q<=24'b110111000001000001001010;
	8'h0x87: q<=24'b110111000001000001001010;
	8'h0x88: q<=24'b110111000001000001001010;
	8'h0x89: q<=24'b110111000001000001001010;
	8'h0x8a: q<=24'b110111000001000001001010;
	8'h0x8b: q<=24'b110111000001000001001010;
	8'h0x8c: q<=24'b110111000001000001001010;
	8'h0x8d: q<=24'b110111000001000001001010;
	8'h0x8e: q<=24'b110111000001000001001010;
	8'h0x8f: q<=24'b110111000001000001001010;
	8'h0x90: q<=24'b110111000001000001001010;
	8'h0x91: q<=24'b110111000001000001001010;
	8'h0x92: q<=24'b110111000001000001001010;
	8'h0x93: q<=24'b110111000001000001001010;
	8'h0x94: q<=24'b000010010010000000110000;
	8'h0x95: q<=24'b000011011100000000110000;
	8'h0x96: q<=24'b100110100000000010010000;
	8'h0x97: q<=24'b000001010011000000001100;
	8'h0x98: q<=24'b000000000010001000000001;
	8'h0x99: q<=24'b000011010011001000110001;
	8'h0x9a: q<=24'b100010000001001001000001;
	8'h0x9b: q<=24'b110110000001000001001010;
	8'h0x9c: q<=24'b110110000001000001001010;
	8'h0x9d: q<=24'b110110000001000001001010;
	8'h0x9e: q<=24'b110110000001000001001010;
	8'h0x9f: q<=24'b110110000001000001001010;
	8'h0xa0: q<=24'b110110000001000001001010;
	8'h0xa1: q<=24'b110110000001000001001010;
	8'h0xa2: q<=24'b110110000001000001001010;
	8'h0xa3: q<=24'b110110000001000001001010;
	8'h0xa4: q<=24'b110110000001000001001010;
	8'h0xa5: q<=24'b110110000001000001001010;
	8'h0xa6: q<=24'b110110000001000001001010;
	8'h0xa7: q<=24'b110110000001000001001010;
	8'h0xa8: q<=24'b110110000001000001001010;
	8'h0xa9: q<=24'b110110000001000001001010;
	8'h0xaa: q<=24'b110110000001000001001010;
	8'h0xab: q<=24'b110010000001000000110000;
	8'h0xac: q<=24'b000010010011000001010000;
	8'h0xad: q<=24'b000011000010000001010000;
	8'h0xae: q<=24'b110010010001000000110000;
	8'h0xaf: q<=24'b101100100010010010000000;
	8'h0xb0: q<=24'b000010010011000001101100;
	8'h0xb1: q<=24'b000010000011000000110001;
	8'h0xb2: q<=24'b101101010000000010010000;
	8'h0xb3: q<=24'b000011110011000000011100;
	8'h0xb4: q<=24'b000010000011100000110000;
	8'h0xb5: q<=24'b001110000001000000110000;
	8'h0xb6: q<=24'b000000000001011100000000;
	8'h0xb7: q<=24'b100110010100010000110000;
	8'h0xb8: q<=24'b100111001100000000110000;
	8'h0xb9: q<=24'b000010000011000000000000;
	8'h0xba: q<=24'b101111110000000010010100;
	8'h0xbb: q<=24'b000000000010000100000000;
	8'h0xbc: q<=24'b011001101000110000110000;
	8'h0xbd: q<=24'b101011001100000000110000;
	8'h0xbe: q<=24'b000010110011000000000000;
	8'h0xbf: q<=24'b011111100000011000110000;
	8'h0xc0: q<=24'b110010000000000010010000;
	8'h0xc1: q<=24'b000011010010000000111100;
	8'h0xc2: q<=24'b000011010010001000110000;
	8'h0xc3: q<=24'b110001110000000010010000;
	8'h0xc4: q<=24'b000011000011001000001100;
	8'h0xc5: q<=24'b110001110010000010011101;
	8'h0xc6: q<=24'b000011010011000000110001;
	8'h0xc7: q<=24'b110010010010000010000101;
	8'h0xc8: q<=24'b000011000011000000000000;
	8'h0xc9: q<=24'b110011000000000010010000;
	8'h0xca: q<=24'b011111001100000000111100;
	8'h0xcb: q<=24'b011111001100001000110001;
	8'h0xcc: q<=24'b011011111100001100110000;
	8'h0xcd: q<=24'b110011010001000100110001;
	8'h0xce: q<=24'b110100101100000010011100;
	8'h0xcf: q<=24'b110011010001000011100000;
	8'h0xd0: q<=24'b000011110011000100111100;
	8'h0xd1: q<=24'b110101010000000010010100;
	8'h0xd2: q<=24'b000011010011000001100000;
	8'h0xd3: q<=24'b110011010010000010000001;
	8'h0xd4: q<=24'b000011110011000100111100;
	8'h0xd5: q<=24'b110110000000000010010000;
	8'h0xd6: q<=24'b000011100011000000011100;
	8'h0xd7: q<=24'b000000000010101000000001;
	8'h0xd8: q<=24'b000000000010100000010000;
	8'h0xd9: q<=24'b000001011011001100110000;
	8'h0xda: q<=24'b000001110011000000000000;
	8'h0xdb: q<=24'b010011100000000001011000;
	8'h0xdc: q<=24'b000010000011000000000000;
	8'h0xdd: q<=24'b010111110000000001011000;
	8'h0xde: q<=24'b111010000000000010010000;
	8'h0xdf: q<=24'b101111100001001000011101;
	8'h0xe0: q<=24'b111111100001001000011101;
	8'h0xe1: q<=24'b111011110001000000000000;
	8'h0xe2: q<=24'b000000000010001000011101;
	8'h0xe3: q<=24'b111001111100000000110000;
	8'h0xe4: q<=24'b111110001100000000110000;
	8'h0xe5: q<=24'b110110100000000010010000;
	8'h0xe6: q<=24'b000001100011000100111100;
	8'h0xe7: q<=24'b000010000011100000010000;
	8'h0xe8: q<=24'b111001001100000000110000;
	8'h0xe9: q<=24'b111101011100000000110000;
	8'h0xea: q<=24'b111001010000000010010100;
	8'h0xeb: q<=24'b000000111011001100110000;
	8'h0xec: q<=24'b111100000000000010010000;
	8'h0xed: q<=24'b000000100001000100110001;
	8'h0xee: q<=24'b000000100011000000011100;
	8'h0xef: q<=24'b000000100011001000110001;
	8'h0xf0: q<=24'b111101000000000010010000;
	8'h0xf1: q<=24'b000100110001000100110001;
	8'h0xf2: q<=24'b000000110011000000011100;
	8'h0xf3: q<=24'b000000110011001000110001;
	8'h0xf4: q<=24'b001011001100000000110000;
	8'h0xf5: q<=24'b001111011100000000110000;
	8'h0xf6: q<=24'b111110100000000010010000;
	8'h0xf7: q<=24'b001000110001000100011101;
	8'h0xf8: q<=24'b001111001100000000110000;
	8'h0xf9: q<=24'b001011011100000000110000;
	8'h0xfa: q<=24'b000011000011000001010000;
	8'h0xfb: q<=24'b000011000011000001010000;
	8'h0xfc: q<=24'b110011010001000000110000;
	8'h0xfd: q<=24'b000011000011000001010000;
	8'h0xfe: q<=24'b110011010001100000110000;
	8'h0xff: q<=24'b000000000000000000000000;
endcase
end
assign dout=q;
endmodule
